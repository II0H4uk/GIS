* SPICE NETLIST
***************************************

.SUBCKT pmos_a_CDNS_5887047866540 1 2 3
** N=3 EP=3 IP=0 FDC=1
M0 2 3 1 1 pmos_a L=2.4e-07 W=1.2e-06 AD=7.2e-13 AS=1.26e-13 PD=1.8e-06 PS=9e-07 w_cont=6e-07 nfing=1 mmm=1 $X=620 $Y=200 $D=5
.ENDS
***************************************
.SUBCKT nmos_a_CDNS_5887047866517
** N=3 EP=0 IP=0 FDC=0
*.SEEDPROM
.ENDS
***************************************
.SUBCKT dn_CDNS_587555745026
** N=2 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT ICV_1
** N=3 EP=0 IP=4 FDC=0
.ENDS
***************************************
.SUBCKT ICV_2
** N=3 EP=0 IP=7 FDC=0
.ENDS
***************************************
.SUBCKT ICV_3
** N=3 EP=0 IP=6 FDC=0
.ENDS
***************************************
.SUBCKT cpoly_n_CDNS_588704786651 1 2
** N=2 EP=2 IP=0 FDC=39
M0 1 2 1 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=1.67141e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=620 $Y=200 $D=22
M1 1 2 1 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=3140 $Y=200 $D=22
M2 1 2 1 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=5660 $Y=200 $D=22
M3 1 2 1 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=8180 $Y=200 $D=22
M4 1 2 1 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=10700 $Y=200 $D=22
M5 1 2 1 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=13220 $Y=200 $D=22
M6 1 2 1 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=15740 $Y=200 $D=22
M7 1 2 1 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=18260 $Y=200 $D=22
M8 1 2 1 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=20780 $Y=200 $D=22
M9 1 2 1 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=23300 $Y=200 $D=22
M10 1 2 1 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=25820 $Y=200 $D=22
M11 1 2 1 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=28340 $Y=200 $D=22
M12 1 2 1 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=30860 $Y=200 $D=22
M13 1 2 1 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=33380 $Y=200 $D=22
M14 1 2 1 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=35900 $Y=200 $D=22
M15 1 2 1 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=38420 $Y=200 $D=22
M16 1 2 1 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=40940 $Y=200 $D=22
M17 1 2 1 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=43460 $Y=200 $D=22
M18 1 2 1 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=45980 $Y=200 $D=22
M19 1 2 1 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=48500 $Y=200 $D=22
M20 1 2 1 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=51020 $Y=200 $D=22
M21 1 2 1 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=53540 $Y=200 $D=22
M22 1 2 1 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=56060 $Y=200 $D=22
M23 1 2 1 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=58580 $Y=200 $D=22
M24 1 2 1 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=61100 $Y=200 $D=22
M25 1 2 1 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=63620 $Y=200 $D=22
M26 1 2 1 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=66140 $Y=200 $D=22
M27 1 2 1 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=68660 $Y=200 $D=22
M28 1 2 1 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=71180 $Y=200 $D=22
M29 1 2 1 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=73700 $Y=200 $D=22
M30 1 2 1 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=76220 $Y=200 $D=22
M31 1 2 1 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=78740 $Y=200 $D=22
M32 1 2 1 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=81260 $Y=200 $D=22
M33 1 2 1 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=83780 $Y=200 $D=22
M34 1 2 1 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=86300 $Y=200 $D=22
M35 1 2 1 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=88820 $Y=200 $D=22
M36 1 2 1 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=91340 $Y=200 $D=22
M37 1 2 1 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=93860 $Y=200 $D=22
M38 1 2 1 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=2.304e-12 ps=2.88e-06 pd=5.14246e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=96380 $Y=200 $D=22
.ENDS
***************************************
.SUBCKT cpoly_p_CDNS_588704786650 1 2
** N=2 EP=2 IP=0 FDC=39
M0 1 2 1 cpoly_p w=8.62e-06 l=2e-06 c=1.08536e-13 as=1.21314e-13 ad=7.488e-13 ps=1.44e-06 pd=1.21456e-06 sim_w=2.88e-06 m_per_maxw=2.99306 numb_sub_cont=4 nfing=1 $X=620 $Y=200 $D=21
M1 1 2 1 cpoly_p w=8.62e-06 l=2e-06 c=1.08536e-13 as=1.53388e-13 ad=7.488e-13 ps=1.44e-06 pd=1.21456e-06 sim_w=2.88e-06 m_per_maxw=2.99306 numb_sub_cont=4 nfing=1 $X=3140 $Y=200 $D=21
M2 1 2 1 cpoly_p w=8.62e-06 l=2e-06 c=1.08536e-13 as=1.53388e-13 ad=7.488e-13 ps=1.44e-06 pd=1.21456e-06 sim_w=2.88e-06 m_per_maxw=2.99306 numb_sub_cont=4 nfing=1 $X=5660 $Y=200 $D=21
M3 1 2 1 cpoly_p w=8.62e-06 l=2e-06 c=1.08536e-13 as=1.53388e-13 ad=7.488e-13 ps=1.44e-06 pd=1.21456e-06 sim_w=2.88e-06 m_per_maxw=2.99306 numb_sub_cont=4 nfing=1 $X=8180 $Y=200 $D=21
M4 1 2 1 cpoly_p w=8.62e-06 l=2e-06 c=1.08536e-13 as=1.53388e-13 ad=7.488e-13 ps=1.44e-06 pd=1.21456e-06 sim_w=2.88e-06 m_per_maxw=2.99306 numb_sub_cont=4 nfing=1 $X=10700 $Y=200 $D=21
M5 1 2 1 cpoly_p w=8.62e-06 l=2e-06 c=1.08536e-13 as=1.53388e-13 ad=7.488e-13 ps=1.44e-06 pd=1.21456e-06 sim_w=2.88e-06 m_per_maxw=2.99306 numb_sub_cont=4 nfing=1 $X=13220 $Y=200 $D=21
M6 1 2 1 cpoly_p w=8.62e-06 l=2e-06 c=1.08536e-13 as=1.53388e-13 ad=7.488e-13 ps=1.44e-06 pd=1.21456e-06 sim_w=2.88e-06 m_per_maxw=2.99306 numb_sub_cont=4 nfing=1 $X=15740 $Y=200 $D=21
M7 1 2 1 cpoly_p w=8.62e-06 l=2e-06 c=1.08536e-13 as=1.53388e-13 ad=7.488e-13 ps=1.44e-06 pd=1.21456e-06 sim_w=2.88e-06 m_per_maxw=2.99306 numb_sub_cont=4 nfing=1 $X=18260 $Y=200 $D=21
M8 1 2 1 cpoly_p w=8.62e-06 l=2e-06 c=1.08536e-13 as=1.53388e-13 ad=7.488e-13 ps=1.44e-06 pd=1.21456e-06 sim_w=2.88e-06 m_per_maxw=2.99306 numb_sub_cont=4 nfing=1 $X=20780 $Y=200 $D=21
M9 1 2 1 cpoly_p w=8.62e-06 l=2e-06 c=1.08536e-13 as=1.53388e-13 ad=7.488e-13 ps=1.44e-06 pd=1.21456e-06 sim_w=2.88e-06 m_per_maxw=2.99306 numb_sub_cont=4 nfing=1 $X=23300 $Y=200 $D=21
M10 1 2 1 cpoly_p w=8.62e-06 l=2e-06 c=1.08536e-13 as=1.53388e-13 ad=7.488e-13 ps=1.44e-06 pd=1.21456e-06 sim_w=2.88e-06 m_per_maxw=2.99306 numb_sub_cont=4 nfing=1 $X=25820 $Y=200 $D=21
M11 1 2 1 cpoly_p w=8.62e-06 l=2e-06 c=1.08536e-13 as=1.53388e-13 ad=7.488e-13 ps=1.44e-06 pd=1.21456e-06 sim_w=2.88e-06 m_per_maxw=2.99306 numb_sub_cont=4 nfing=1 $X=28340 $Y=200 $D=21
M12 1 2 1 cpoly_p w=8.62e-06 l=2e-06 c=1.08536e-13 as=1.53388e-13 ad=7.488e-13 ps=1.44e-06 pd=1.21456e-06 sim_w=2.88e-06 m_per_maxw=2.99306 numb_sub_cont=4 nfing=1 $X=30860 $Y=200 $D=21
M13 1 2 1 cpoly_p w=8.62e-06 l=2e-06 c=1.08536e-13 as=1.53388e-13 ad=7.488e-13 ps=1.44e-06 pd=1.21456e-06 sim_w=2.88e-06 m_per_maxw=2.99306 numb_sub_cont=4 nfing=1 $X=33380 $Y=200 $D=21
M14 1 2 1 cpoly_p w=8.62e-06 l=2e-06 c=1.08536e-13 as=1.53388e-13 ad=7.488e-13 ps=1.44e-06 pd=1.21456e-06 sim_w=2.88e-06 m_per_maxw=2.99306 numb_sub_cont=4 nfing=1 $X=35900 $Y=200 $D=21
M15 1 2 1 cpoly_p w=8.62e-06 l=2e-06 c=1.08536e-13 as=1.53388e-13 ad=7.488e-13 ps=1.44e-06 pd=1.21456e-06 sim_w=2.88e-06 m_per_maxw=2.99306 numb_sub_cont=4 nfing=1 $X=38420 $Y=200 $D=21
M16 1 2 1 cpoly_p w=8.62e-06 l=2e-06 c=1.08536e-13 as=1.53388e-13 ad=7.488e-13 ps=1.44e-06 pd=1.21456e-06 sim_w=2.88e-06 m_per_maxw=2.99306 numb_sub_cont=4 nfing=1 $X=40940 $Y=200 $D=21
M17 1 2 1 cpoly_p w=8.62e-06 l=2e-06 c=1.08536e-13 as=1.53388e-13 ad=7.488e-13 ps=1.44e-06 pd=1.21456e-06 sim_w=2.88e-06 m_per_maxw=2.99306 numb_sub_cont=4 nfing=1 $X=43460 $Y=200 $D=21
M18 1 2 1 cpoly_p w=8.62e-06 l=2e-06 c=1.08536e-13 as=1.53388e-13 ad=7.488e-13 ps=1.44e-06 pd=1.21456e-06 sim_w=2.88e-06 m_per_maxw=2.99306 numb_sub_cont=4 nfing=1 $X=45980 $Y=200 $D=21
M19 1 2 1 cpoly_p w=8.62e-06 l=2e-06 c=1.08536e-13 as=1.53388e-13 ad=7.488e-13 ps=1.44e-06 pd=1.21456e-06 sim_w=2.88e-06 m_per_maxw=2.99306 numb_sub_cont=4 nfing=1 $X=48500 $Y=200 $D=21
M20 1 2 1 cpoly_p w=8.62e-06 l=2e-06 c=1.08536e-13 as=1.53388e-13 ad=7.488e-13 ps=1.44e-06 pd=1.21456e-06 sim_w=2.88e-06 m_per_maxw=2.99306 numb_sub_cont=4 nfing=1 $X=51020 $Y=200 $D=21
M21 1 2 1 cpoly_p w=8.62e-06 l=2e-06 c=1.08536e-13 as=1.53388e-13 ad=7.488e-13 ps=1.44e-06 pd=1.21456e-06 sim_w=2.88e-06 m_per_maxw=2.99306 numb_sub_cont=4 nfing=1 $X=53540 $Y=200 $D=21
M22 1 2 1 cpoly_p w=8.62e-06 l=2e-06 c=1.08536e-13 as=1.53388e-13 ad=7.488e-13 ps=1.44e-06 pd=1.21456e-06 sim_w=2.88e-06 m_per_maxw=2.99306 numb_sub_cont=4 nfing=1 $X=56060 $Y=200 $D=21
M23 1 2 1 cpoly_p w=8.62e-06 l=2e-06 c=1.08536e-13 as=1.53388e-13 ad=7.488e-13 ps=1.44e-06 pd=1.21456e-06 sim_w=2.88e-06 m_per_maxw=2.99306 numb_sub_cont=4 nfing=1 $X=58580 $Y=200 $D=21
M24 1 2 1 cpoly_p w=8.62e-06 l=2e-06 c=1.08536e-13 as=1.53388e-13 ad=7.488e-13 ps=1.44e-06 pd=1.21456e-06 sim_w=2.88e-06 m_per_maxw=2.99306 numb_sub_cont=4 nfing=1 $X=61100 $Y=200 $D=21
M25 1 2 1 cpoly_p w=8.62e-06 l=2e-06 c=1.08536e-13 as=1.53388e-13 ad=7.488e-13 ps=1.44e-06 pd=1.21456e-06 sim_w=2.88e-06 m_per_maxw=2.99306 numb_sub_cont=4 nfing=1 $X=63620 $Y=200 $D=21
M26 1 2 1 cpoly_p w=8.62e-06 l=2e-06 c=1.08536e-13 as=1.53388e-13 ad=7.488e-13 ps=1.44e-06 pd=1.21456e-06 sim_w=2.88e-06 m_per_maxw=2.99306 numb_sub_cont=4 nfing=1 $X=66140 $Y=200 $D=21
M27 1 2 1 cpoly_p w=8.62e-06 l=2e-06 c=1.08536e-13 as=1.53388e-13 ad=7.488e-13 ps=1.44e-06 pd=1.21456e-06 sim_w=2.88e-06 m_per_maxw=2.99306 numb_sub_cont=4 nfing=1 $X=68660 $Y=200 $D=21
M28 1 2 1 cpoly_p w=8.62e-06 l=2e-06 c=1.08536e-13 as=1.53388e-13 ad=7.488e-13 ps=1.44e-06 pd=1.21456e-06 sim_w=2.88e-06 m_per_maxw=2.99306 numb_sub_cont=4 nfing=1 $X=71180 $Y=200 $D=21
M29 1 2 1 cpoly_p w=8.62e-06 l=2e-06 c=1.08536e-13 as=1.53388e-13 ad=7.488e-13 ps=1.44e-06 pd=1.21456e-06 sim_w=2.88e-06 m_per_maxw=2.99306 numb_sub_cont=4 nfing=1 $X=73700 $Y=200 $D=21
M30 1 2 1 cpoly_p w=8.62e-06 l=2e-06 c=1.08536e-13 as=1.53388e-13 ad=7.488e-13 ps=1.44e-06 pd=1.21456e-06 sim_w=2.88e-06 m_per_maxw=2.99306 numb_sub_cont=4 nfing=1 $X=76220 $Y=200 $D=21
M31 1 2 1 cpoly_p w=8.62e-06 l=2e-06 c=1.08536e-13 as=1.53388e-13 ad=7.488e-13 ps=1.44e-06 pd=1.21456e-06 sim_w=2.88e-06 m_per_maxw=2.99306 numb_sub_cont=4 nfing=1 $X=78740 $Y=200 $D=21
M32 1 2 1 cpoly_p w=8.62e-06 l=2e-06 c=1.08536e-13 as=1.53388e-13 ad=7.488e-13 ps=1.44e-06 pd=1.21456e-06 sim_w=2.88e-06 m_per_maxw=2.99306 numb_sub_cont=4 nfing=1 $X=81260 $Y=200 $D=21
M33 1 2 1 cpoly_p w=8.62e-06 l=2e-06 c=1.08536e-13 as=1.53388e-13 ad=7.488e-13 ps=1.44e-06 pd=1.21456e-06 sim_w=2.88e-06 m_per_maxw=2.99306 numb_sub_cont=4 nfing=1 $X=83780 $Y=200 $D=21
M34 1 2 1 cpoly_p w=8.62e-06 l=2e-06 c=1.08536e-13 as=1.53388e-13 ad=7.488e-13 ps=1.44e-06 pd=1.21456e-06 sim_w=2.88e-06 m_per_maxw=2.99306 numb_sub_cont=4 nfing=1 $X=86300 $Y=200 $D=21
M35 1 2 1 cpoly_p w=8.62e-06 l=2e-06 c=1.08536e-13 as=1.53388e-13 ad=7.488e-13 ps=1.44e-06 pd=1.21456e-06 sim_w=2.88e-06 m_per_maxw=2.99306 numb_sub_cont=4 nfing=1 $X=88820 $Y=200 $D=21
M36 1 2 1 cpoly_p w=8.62e-06 l=2e-06 c=1.08536e-13 as=1.53388e-13 ad=7.488e-13 ps=1.44e-06 pd=1.21456e-06 sim_w=2.88e-06 m_per_maxw=2.99306 numb_sub_cont=4 nfing=1 $X=91340 $Y=200 $D=21
M37 1 2 1 cpoly_p w=8.62e-06 l=2e-06 c=1.08536e-13 as=1.53388e-13 ad=7.488e-13 ps=1.44e-06 pd=1.21456e-06 sim_w=2.88e-06 m_per_maxw=2.99306 numb_sub_cont=4 nfing=1 $X=93860 $Y=200 $D=21
M38 1 2 1 cpoly_p w=8.62e-06 l=2e-06 c=1.08536e-13 as=1.53388e-13 ad=1.152e-12 ps=1.44e-06 pd=2.42912e-06 sim_w=2.88e-06 m_per_maxw=2.99306 numb_sub_cont=4 nfing=1 $X=96380 $Y=200 $D=21
.ENDS
***************************************
.SUBCKT VDD_PAD gnd! vdd!
** N=8 EP=2 IP=26 FDC=78
*.CALIBRE ISOLATED NETS: VDD_PAD GND_PAD
X8 vdd! gnd! cpoly_n_CDNS_588704786651 $T=520 333340 0 0 $X=520 $Y=333340
X9 gnd! vdd! cpoly_p_CDNS_588704786650 $T=520 320500 0 0 $X=520 $Y=320500
.ENDS
***************************************
.SUBCKT pmos_a_CDNS_5887047866567
** N=3 EP=0 IP=0 FDC=0
*.SEEDPROM
.ENDS
***************************************
.SUBCKT nmos_a_CDNS_5887047866553 1 2 3
** N=3 EP=3 IP=0 FDC=1
M0 2 3 1 1 nmos_a L=2.4e-07 W=4.8e-06 AD=1.656e-12 AS=1.92e-12 PD=4.14e-06 PS=2.07e-06 w_cont=2.1e-06 nfing=1 source_num=2 $X=620 $Y=200 $D=1
.ENDS
***************************************
.SUBCKT cpoly_n_CDNS_5887047866516
** N=2 EP=0 IP=0 FDC=0
*.SEEDPROM
.ENDS
***************************************
.SUBCKT pmos_a_CDNS_5887047866519
** N=3 EP=0 IP=0 FDC=0
*.SEEDPROM
.ENDS
***************************************
.SUBCKT nmos_a_CDNS_5887047866525
** N=3 EP=0 IP=0 FDC=0
*.SEEDPROM
.ENDS
***************************************
.SUBCKT pmos_a_CDNS_5887047866513
** N=3 EP=0 IP=0 FDC=0
*.SEEDPROM
.ENDS
***************************************
.SUBCKT nmos_a_CDNS_5887047866526
** N=3 EP=0 IP=0 FDC=0
*.SEEDPROM
.ENDS
***************************************
.SUBCKT nmos_a_CDNS_5887047866524
** N=3 EP=0 IP=0 FDC=0
*.SEEDPROM
.ENDS
***************************************
.SUBCKT pmos_a_CDNS_5887047866518
** N=3 EP=0 IP=0 FDC=0
*.SEEDPROM
.ENDS
***************************************
.SUBCKT cpoly_p_CDNS_5887047866511 1 2
** N=2 EP=2 IP=0 FDC=36
M0 1 2 1 cpoly_p w=6e-06 l=2e-06 c=8.0712e-14 as=1.68e-13 ad=7.488e-13 ps=1.44e-06 pd=1.13684e-06 sim_w=2.88e-06 m_per_maxw=2.08333 numb_sub_cont=4 nfing=1 $X=620 $Y=200 $D=21
M1 1 2 1 cpoly_p w=6e-06 l=2e-06 c=8.0712e-14 as=2.1408e-13 ad=7.488e-13 ps=1.44e-06 pd=1.13684e-06 sim_w=2.88e-06 m_per_maxw=2.08333 numb_sub_cont=4 nfing=1 $X=3140 $Y=200 $D=21
M2 1 2 1 cpoly_p w=6e-06 l=2e-06 c=8.0712e-14 as=2.1408e-13 ad=7.488e-13 ps=1.44e-06 pd=1.13684e-06 sim_w=2.88e-06 m_per_maxw=2.08333 numb_sub_cont=4 nfing=1 $X=5660 $Y=200 $D=21
M3 1 2 1 cpoly_p w=6e-06 l=2e-06 c=8.0712e-14 as=2.1408e-13 ad=7.488e-13 ps=1.44e-06 pd=1.13684e-06 sim_w=2.88e-06 m_per_maxw=2.08333 numb_sub_cont=4 nfing=1 $X=8180 $Y=200 $D=21
M4 1 2 1 cpoly_p w=6e-06 l=2e-06 c=8.0712e-14 as=2.1408e-13 ad=7.488e-13 ps=1.44e-06 pd=1.13684e-06 sim_w=2.88e-06 m_per_maxw=2.08333 numb_sub_cont=4 nfing=1 $X=10700 $Y=200 $D=21
M5 1 2 1 cpoly_p w=6e-06 l=2e-06 c=8.0712e-14 as=2.1408e-13 ad=7.488e-13 ps=1.44e-06 pd=1.13684e-06 sim_w=2.88e-06 m_per_maxw=2.08333 numb_sub_cont=4 nfing=1 $X=13220 $Y=200 $D=21
M6 1 2 1 cpoly_p w=6e-06 l=2e-06 c=8.0712e-14 as=2.1408e-13 ad=7.488e-13 ps=1.44e-06 pd=1.13684e-06 sim_w=2.88e-06 m_per_maxw=2.08333 numb_sub_cont=4 nfing=1 $X=15740 $Y=200 $D=21
M7 1 2 1 cpoly_p w=6e-06 l=2e-06 c=8.0712e-14 as=2.1408e-13 ad=7.488e-13 ps=1.44e-06 pd=1.13684e-06 sim_w=2.88e-06 m_per_maxw=2.08333 numb_sub_cont=4 nfing=1 $X=18260 $Y=200 $D=21
M8 1 2 1 cpoly_p w=6e-06 l=2e-06 c=8.0712e-14 as=2.1408e-13 ad=7.488e-13 ps=1.44e-06 pd=1.13684e-06 sim_w=2.88e-06 m_per_maxw=2.08333 numb_sub_cont=4 nfing=1 $X=20780 $Y=200 $D=21
M9 1 2 1 cpoly_p w=6e-06 l=2e-06 c=8.0712e-14 as=2.1408e-13 ad=7.488e-13 ps=1.44e-06 pd=1.13684e-06 sim_w=2.88e-06 m_per_maxw=2.08333 numb_sub_cont=4 nfing=1 $X=23300 $Y=200 $D=21
M10 1 2 1 cpoly_p w=6e-06 l=2e-06 c=8.0712e-14 as=2.1408e-13 ad=7.488e-13 ps=1.44e-06 pd=1.13684e-06 sim_w=2.88e-06 m_per_maxw=2.08333 numb_sub_cont=4 nfing=1 $X=25820 $Y=200 $D=21
M11 1 2 1 cpoly_p w=6e-06 l=2e-06 c=8.0712e-14 as=2.1408e-13 ad=7.488e-13 ps=1.44e-06 pd=1.13684e-06 sim_w=2.88e-06 m_per_maxw=2.08333 numb_sub_cont=4 nfing=1 $X=28340 $Y=200 $D=21
M12 1 2 1 cpoly_p w=6e-06 l=2e-06 c=8.0712e-14 as=2.1408e-13 ad=7.488e-13 ps=1.44e-06 pd=1.13684e-06 sim_w=2.88e-06 m_per_maxw=2.08333 numb_sub_cont=4 nfing=1 $X=30860 $Y=200 $D=21
M13 1 2 1 cpoly_p w=6e-06 l=2e-06 c=8.0712e-14 as=2.1408e-13 ad=7.488e-13 ps=1.44e-06 pd=1.13684e-06 sim_w=2.88e-06 m_per_maxw=2.08333 numb_sub_cont=4 nfing=1 $X=33380 $Y=200 $D=21
M14 1 2 1 cpoly_p w=6e-06 l=2e-06 c=8.0712e-14 as=2.1408e-13 ad=7.488e-13 ps=1.44e-06 pd=1.13684e-06 sim_w=2.88e-06 m_per_maxw=2.08333 numb_sub_cont=4 nfing=1 $X=35900 $Y=200 $D=21
M15 1 2 1 cpoly_p w=6e-06 l=2e-06 c=8.0712e-14 as=2.1408e-13 ad=7.488e-13 ps=1.44e-06 pd=1.13684e-06 sim_w=2.88e-06 m_per_maxw=2.08333 numb_sub_cont=4 nfing=1 $X=38420 $Y=200 $D=21
M16 1 2 1 cpoly_p w=6e-06 l=2e-06 c=8.0712e-14 as=2.1408e-13 ad=7.488e-13 ps=1.44e-06 pd=1.13684e-06 sim_w=2.88e-06 m_per_maxw=2.08333 numb_sub_cont=4 nfing=1 $X=40940 $Y=200 $D=21
M17 1 2 1 cpoly_p w=6e-06 l=2e-06 c=8.0712e-14 as=2.1408e-13 ad=7.488e-13 ps=1.44e-06 pd=1.13684e-06 sim_w=2.88e-06 m_per_maxw=2.08333 numb_sub_cont=4 nfing=1 $X=43460 $Y=200 $D=21
M18 1 2 1 cpoly_p w=6e-06 l=2e-06 c=8.0712e-14 as=2.1408e-13 ad=7.488e-13 ps=1.44e-06 pd=1.13684e-06 sim_w=2.88e-06 m_per_maxw=2.08333 numb_sub_cont=4 nfing=1 $X=45980 $Y=200 $D=21
M19 1 2 1 cpoly_p w=6e-06 l=2e-06 c=8.0712e-14 as=2.1408e-13 ad=7.488e-13 ps=1.44e-06 pd=1.13684e-06 sim_w=2.88e-06 m_per_maxw=2.08333 numb_sub_cont=4 nfing=1 $X=48500 $Y=200 $D=21
M20 1 2 1 cpoly_p w=6e-06 l=2e-06 c=8.0712e-14 as=2.1408e-13 ad=7.488e-13 ps=1.44e-06 pd=1.13684e-06 sim_w=2.88e-06 m_per_maxw=2.08333 numb_sub_cont=4 nfing=1 $X=51020 $Y=200 $D=21
M21 1 2 1 cpoly_p w=6e-06 l=2e-06 c=8.0712e-14 as=2.1408e-13 ad=7.488e-13 ps=1.44e-06 pd=1.13684e-06 sim_w=2.88e-06 m_per_maxw=2.08333 numb_sub_cont=4 nfing=1 $X=53540 $Y=200 $D=21
M22 1 2 1 cpoly_p w=6e-06 l=2e-06 c=8.0712e-14 as=2.1408e-13 ad=7.488e-13 ps=1.44e-06 pd=1.13684e-06 sim_w=2.88e-06 m_per_maxw=2.08333 numb_sub_cont=4 nfing=1 $X=56060 $Y=200 $D=21
M23 1 2 1 cpoly_p w=6e-06 l=2e-06 c=8.0712e-14 as=2.1408e-13 ad=7.488e-13 ps=1.44e-06 pd=1.13684e-06 sim_w=2.88e-06 m_per_maxw=2.08333 numb_sub_cont=4 nfing=1 $X=58580 $Y=200 $D=21
M24 1 2 1 cpoly_p w=6e-06 l=2e-06 c=8.0712e-14 as=2.1408e-13 ad=7.488e-13 ps=1.44e-06 pd=1.13684e-06 sim_w=2.88e-06 m_per_maxw=2.08333 numb_sub_cont=4 nfing=1 $X=61100 $Y=200 $D=21
M25 1 2 1 cpoly_p w=6e-06 l=2e-06 c=8.0712e-14 as=2.1408e-13 ad=7.488e-13 ps=1.44e-06 pd=1.13684e-06 sim_w=2.88e-06 m_per_maxw=2.08333 numb_sub_cont=4 nfing=1 $X=63620 $Y=200 $D=21
M26 1 2 1 cpoly_p w=6e-06 l=2e-06 c=8.0712e-14 as=2.1408e-13 ad=7.488e-13 ps=1.44e-06 pd=1.13684e-06 sim_w=2.88e-06 m_per_maxw=2.08333 numb_sub_cont=4 nfing=1 $X=66140 $Y=200 $D=21
M27 1 2 1 cpoly_p w=6e-06 l=2e-06 c=8.0712e-14 as=2.1408e-13 ad=7.488e-13 ps=1.44e-06 pd=1.13684e-06 sim_w=2.88e-06 m_per_maxw=2.08333 numb_sub_cont=4 nfing=1 $X=68660 $Y=200 $D=21
M28 1 2 1 cpoly_p w=6e-06 l=2e-06 c=8.0712e-14 as=2.1408e-13 ad=7.488e-13 ps=1.44e-06 pd=1.13684e-06 sim_w=2.88e-06 m_per_maxw=2.08333 numb_sub_cont=4 nfing=1 $X=71180 $Y=200 $D=21
M29 1 2 1 cpoly_p w=6e-06 l=2e-06 c=8.0712e-14 as=2.1408e-13 ad=7.488e-13 ps=1.44e-06 pd=1.13684e-06 sim_w=2.88e-06 m_per_maxw=2.08333 numb_sub_cont=4 nfing=1 $X=73700 $Y=200 $D=21
M30 1 2 1 cpoly_p w=6e-06 l=2e-06 c=8.0712e-14 as=2.1408e-13 ad=7.488e-13 ps=1.44e-06 pd=1.13684e-06 sim_w=2.88e-06 m_per_maxw=2.08333 numb_sub_cont=4 nfing=1 $X=76220 $Y=200 $D=21
M31 1 2 1 cpoly_p w=6e-06 l=2e-06 c=8.0712e-14 as=2.1408e-13 ad=7.488e-13 ps=1.44e-06 pd=1.13684e-06 sim_w=2.88e-06 m_per_maxw=2.08333 numb_sub_cont=4 nfing=1 $X=78740 $Y=200 $D=21
M32 1 2 1 cpoly_p w=6e-06 l=2e-06 c=8.0712e-14 as=2.1408e-13 ad=7.488e-13 ps=1.44e-06 pd=1.13684e-06 sim_w=2.88e-06 m_per_maxw=2.08333 numb_sub_cont=4 nfing=1 $X=81260 $Y=200 $D=21
M33 1 2 1 cpoly_p w=6e-06 l=2e-06 c=8.0712e-14 as=2.1408e-13 ad=7.488e-13 ps=1.44e-06 pd=1.13684e-06 sim_w=2.88e-06 m_per_maxw=2.08333 numb_sub_cont=4 nfing=1 $X=83780 $Y=200 $D=21
M34 1 2 1 cpoly_p w=6e-06 l=2e-06 c=8.0712e-14 as=2.1408e-13 ad=7.488e-13 ps=1.44e-06 pd=1.13684e-06 sim_w=2.88e-06 m_per_maxw=2.08333 numb_sub_cont=4 nfing=1 $X=86300 $Y=200 $D=21
M35 1 2 1 cpoly_p w=6e-06 l=2e-06 c=8.0712e-14 as=1.68e-13 ad=7.488e-13 ps=1.44e-06 pd=1.13684e-06 sim_w=2.88e-06 m_per_maxw=2.08333 numb_sub_cont=4 nfing=1 $X=88820 $Y=200 $D=21
.ENDS
***************************************
.SUBCKT cpoly_n_CDNS_5887047866514 1 2
** N=2 EP=2 IP=0 FDC=39
M0 1 2 1 cpoly_n w=6e-06 l=2e-06 c=7.5402e-14 as=2.4e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.4338e-06 sim_w=5.76e-06 m_per_maxw=1.04167 numb_sub_cont=3 nfing=1 $X=620 $Y=200 $D=22
M1 1 2 1 cpoly_n w=6e-06 l=2e-06 c=7.5402e-14 as=3.0336e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.4338e-06 sim_w=5.76e-06 m_per_maxw=1.04167 numb_sub_cont=3 nfing=1 $X=3140 $Y=200 $D=22
M2 1 2 1 cpoly_n w=6e-06 l=2e-06 c=7.5402e-14 as=3.0336e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.4338e-06 sim_w=5.76e-06 m_per_maxw=1.04167 numb_sub_cont=3 nfing=1 $X=5660 $Y=200 $D=22
M3 1 2 1 cpoly_n w=6e-06 l=2e-06 c=7.5402e-14 as=3.0336e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.4338e-06 sim_w=5.76e-06 m_per_maxw=1.04167 numb_sub_cont=3 nfing=1 $X=8180 $Y=200 $D=22
M4 1 2 1 cpoly_n w=6e-06 l=2e-06 c=7.5402e-14 as=3.0336e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.4338e-06 sim_w=5.76e-06 m_per_maxw=1.04167 numb_sub_cont=3 nfing=1 $X=10700 $Y=200 $D=22
M5 1 2 1 cpoly_n w=6e-06 l=2e-06 c=7.5402e-14 as=3.0336e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.4338e-06 sim_w=5.76e-06 m_per_maxw=1.04167 numb_sub_cont=3 nfing=1 $X=13220 $Y=200 $D=22
M6 1 2 1 cpoly_n w=6e-06 l=2e-06 c=7.5402e-14 as=3.0336e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.4338e-06 sim_w=5.76e-06 m_per_maxw=1.04167 numb_sub_cont=3 nfing=1 $X=15740 $Y=200 $D=22
M7 1 2 1 cpoly_n w=6e-06 l=2e-06 c=7.5402e-14 as=3.0336e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.4338e-06 sim_w=5.76e-06 m_per_maxw=1.04167 numb_sub_cont=3 nfing=1 $X=18260 $Y=200 $D=22
M8 1 2 1 cpoly_n w=6e-06 l=2e-06 c=7.5402e-14 as=3.0336e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.4338e-06 sim_w=5.76e-06 m_per_maxw=1.04167 numb_sub_cont=3 nfing=1 $X=20780 $Y=200 $D=22
M9 1 2 1 cpoly_n w=6e-06 l=2e-06 c=7.5402e-14 as=3.0336e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.4338e-06 sim_w=5.76e-06 m_per_maxw=1.04167 numb_sub_cont=3 nfing=1 $X=23300 $Y=200 $D=22
M10 1 2 1 cpoly_n w=6e-06 l=2e-06 c=7.5402e-14 as=3.0336e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.4338e-06 sim_w=5.76e-06 m_per_maxw=1.04167 numb_sub_cont=3 nfing=1 $X=25820 $Y=200 $D=22
M11 1 2 1 cpoly_n w=6e-06 l=2e-06 c=7.5402e-14 as=3.0336e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.4338e-06 sim_w=5.76e-06 m_per_maxw=1.04167 numb_sub_cont=3 nfing=1 $X=28340 $Y=200 $D=22
M12 1 2 1 cpoly_n w=6e-06 l=2e-06 c=7.5402e-14 as=3.0336e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.4338e-06 sim_w=5.76e-06 m_per_maxw=1.04167 numb_sub_cont=3 nfing=1 $X=30860 $Y=200 $D=22
M13 1 2 1 cpoly_n w=6e-06 l=2e-06 c=7.5402e-14 as=3.0336e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.4338e-06 sim_w=5.76e-06 m_per_maxw=1.04167 numb_sub_cont=3 nfing=1 $X=33380 $Y=200 $D=22
M14 1 2 1 cpoly_n w=6e-06 l=2e-06 c=7.5402e-14 as=3.0336e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.4338e-06 sim_w=5.76e-06 m_per_maxw=1.04167 numb_sub_cont=3 nfing=1 $X=35900 $Y=200 $D=22
M15 1 2 1 cpoly_n w=6e-06 l=2e-06 c=7.5402e-14 as=3.0336e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.4338e-06 sim_w=5.76e-06 m_per_maxw=1.04167 numb_sub_cont=3 nfing=1 $X=38420 $Y=200 $D=22
M16 1 2 1 cpoly_n w=6e-06 l=2e-06 c=7.5402e-14 as=3.0336e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.4338e-06 sim_w=5.76e-06 m_per_maxw=1.04167 numb_sub_cont=3 nfing=1 $X=40940 $Y=200 $D=22
M17 1 2 1 cpoly_n w=6e-06 l=2e-06 c=7.5402e-14 as=3.0336e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.4338e-06 sim_w=5.76e-06 m_per_maxw=1.04167 numb_sub_cont=3 nfing=1 $X=43460 $Y=200 $D=22
M18 1 2 1 cpoly_n w=6e-06 l=2e-06 c=7.5402e-14 as=3.0336e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.4338e-06 sim_w=5.76e-06 m_per_maxw=1.04167 numb_sub_cont=3 nfing=1 $X=45980 $Y=200 $D=22
M19 1 2 1 cpoly_n w=6e-06 l=2e-06 c=7.5402e-14 as=3.0336e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.4338e-06 sim_w=5.76e-06 m_per_maxw=1.04167 numb_sub_cont=3 nfing=1 $X=48500 $Y=200 $D=22
M20 1 2 1 cpoly_n w=6e-06 l=2e-06 c=7.5402e-14 as=3.0336e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.4338e-06 sim_w=5.76e-06 m_per_maxw=1.04167 numb_sub_cont=3 nfing=1 $X=51020 $Y=200 $D=22
M21 1 2 1 cpoly_n w=6e-06 l=2e-06 c=7.5402e-14 as=3.0336e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.4338e-06 sim_w=5.76e-06 m_per_maxw=1.04167 numb_sub_cont=3 nfing=1 $X=53540 $Y=200 $D=22
M22 1 2 1 cpoly_n w=6e-06 l=2e-06 c=7.5402e-14 as=3.0336e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.4338e-06 sim_w=5.76e-06 m_per_maxw=1.04167 numb_sub_cont=3 nfing=1 $X=56060 $Y=200 $D=22
M23 1 2 1 cpoly_n w=6e-06 l=2e-06 c=7.5402e-14 as=3.0336e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.4338e-06 sim_w=5.76e-06 m_per_maxw=1.04167 numb_sub_cont=3 nfing=1 $X=58580 $Y=200 $D=22
M24 1 2 1 cpoly_n w=6e-06 l=2e-06 c=7.5402e-14 as=3.0336e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.4338e-06 sim_w=5.76e-06 m_per_maxw=1.04167 numb_sub_cont=3 nfing=1 $X=61100 $Y=200 $D=22
M25 1 2 1 cpoly_n w=6e-06 l=2e-06 c=7.5402e-14 as=3.0336e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.4338e-06 sim_w=5.76e-06 m_per_maxw=1.04167 numb_sub_cont=3 nfing=1 $X=63620 $Y=200 $D=22
M26 1 2 1 cpoly_n w=6e-06 l=2e-06 c=7.5402e-14 as=3.0336e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.4338e-06 sim_w=5.76e-06 m_per_maxw=1.04167 numb_sub_cont=3 nfing=1 $X=66140 $Y=200 $D=22
M27 1 2 1 cpoly_n w=6e-06 l=2e-06 c=7.5402e-14 as=3.0336e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.4338e-06 sim_w=5.76e-06 m_per_maxw=1.04167 numb_sub_cont=3 nfing=1 $X=68660 $Y=200 $D=22
M28 1 2 1 cpoly_n w=6e-06 l=2e-06 c=7.5402e-14 as=3.0336e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.4338e-06 sim_w=5.76e-06 m_per_maxw=1.04167 numb_sub_cont=3 nfing=1 $X=71180 $Y=200 $D=22
M29 1 2 1 cpoly_n w=6e-06 l=2e-06 c=7.5402e-14 as=3.0336e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.4338e-06 sim_w=5.76e-06 m_per_maxw=1.04167 numb_sub_cont=3 nfing=1 $X=73700 $Y=200 $D=22
M30 1 2 1 cpoly_n w=6e-06 l=2e-06 c=7.5402e-14 as=3.0336e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.4338e-06 sim_w=5.76e-06 m_per_maxw=1.04167 numb_sub_cont=3 nfing=1 $X=76220 $Y=200 $D=22
M31 1 2 1 cpoly_n w=6e-06 l=2e-06 c=7.5402e-14 as=3.0336e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.4338e-06 sim_w=5.76e-06 m_per_maxw=1.04167 numb_sub_cont=3 nfing=1 $X=78740 $Y=200 $D=22
M32 1 2 1 cpoly_n w=6e-06 l=2e-06 c=7.5402e-14 as=3.0336e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.4338e-06 sim_w=5.76e-06 m_per_maxw=1.04167 numb_sub_cont=3 nfing=1 $X=81260 $Y=200 $D=22
M33 1 2 1 cpoly_n w=6e-06 l=2e-06 c=7.5402e-14 as=3.0336e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.4338e-06 sim_w=5.76e-06 m_per_maxw=1.04167 numb_sub_cont=3 nfing=1 $X=83780 $Y=200 $D=22
M34 1 2 1 cpoly_n w=6e-06 l=2e-06 c=7.5402e-14 as=3.0336e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.4338e-06 sim_w=5.76e-06 m_per_maxw=1.04167 numb_sub_cont=3 nfing=1 $X=86300 $Y=200 $D=22
M35 1 2 1 cpoly_n w=6e-06 l=2e-06 c=7.5402e-14 as=3.0336e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.4338e-06 sim_w=5.76e-06 m_per_maxw=1.04167 numb_sub_cont=3 nfing=1 $X=88820 $Y=200 $D=22
M36 1 2 1 cpoly_n w=6e-06 l=2e-06 c=7.5402e-14 as=3.0336e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.4338e-06 sim_w=5.76e-06 m_per_maxw=1.04167 numb_sub_cont=3 nfing=1 $X=91340 $Y=200 $D=22
M37 1 2 1 cpoly_n w=6e-06 l=2e-06 c=7.5402e-14 as=3.0336e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.4338e-06 sim_w=5.76e-06 m_per_maxw=1.04167 numb_sub_cont=3 nfing=1 $X=93860 $Y=200 $D=22
M38 1 2 1 cpoly_n w=6e-06 l=2e-06 c=7.5402e-14 as=3.0336e-13 ad=2.304e-12 ps=2.88e-06 pd=4.86761e-06 sim_w=5.76e-06 m_per_maxw=1.04167 numb_sub_cont=3 nfing=1 $X=96380 $Y=200 $D=22
.ENDS
***************************************
.SUBCKT dn_CDNS_588704786659
** N=2 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT ICV_4
** N=3 EP=0 IP=4 FDC=0
.ENDS
***************************************
.SUBCKT dn_CDNS_588704786658
** N=2 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT ICV_5
** N=3 EP=0 IP=6 FDC=0
.ENDS
***************************************
.SUBCKT dn_CDNS_5887047866510
** N=2 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT PAD PAD In
** N=10 EP=2 IP=106 FDC=1
*.CALIBRE ISOLATED NETS: gnd1 vdd1 gnd2 vdd2
R0 PAD In 287.224 L=1e-05 W=4e-06 m=1 $[rnpoly] $X=2620 $Y=315480 $D=18
.ENDS
***************************************
.SUBCKT PADIN_WE nATD nClk nWE gnd! vdd! NWR WEN
** N=28 EP=7 IP=163 FDC=217
M0 25 11 gnd! gnd! nmos_a L=2.4e-07 W=2.4e-06 AD=1.4e-12 AS=9.6e-13 PD=3.5e-06 PS=1.75e-06 w_cont=1.1e-06 nfing=1 source_num=2 $X=60860 $Y=327340 $D=1
M1 26 13 25 25 nmos_a L=2.4e-07 W=2.4e-06 AD=1.4e-12 AS=9.6e-13 PD=3.5e-06 PS=1.75e-06 w_cont=1.1e-06 nfing=1 source_num=2 $X=62300 $Y=327340 $D=1
M2 27 12 26 26 nmos_a L=2.4e-07 W=2.4e-06 AD=1.4e-12 AS=9.6e-13 PD=3.5e-06 PS=1.75e-06 w_cont=1.1e-06 nfing=1 source_num=2 $X=63740 $Y=327340 $D=1
M3 nATD 17 gnd! gnd! nmos_a L=2.4e-07 W=1.2e-06 AD=7.2e-13 AS=4.8e-13 PD=1.8e-06 PS=9e-07 w_cont=6e-07 nfing=1 source_num=2 $X=14960 $Y=327320 $D=1
M4 20 8 gnd! gnd! nmos_a L=2.4e-07 W=1.2e-06 AD=7.2e-13 AS=4.8e-13 PD=1.8e-06 PS=9e-07 w_cont=6e-07 nfing=1 source_num=2 $X=27360 $Y=328420 $D=1
M5 21 13 gnd! gnd! nmos_a L=2.4e-07 W=1.2e-06 AD=7.2e-13 AS=4.8e-13 PD=1.8e-06 PS=9e-07 w_cont=6e-07 nfing=1 source_num=2 $X=49760 $Y=328380 $D=1
M6 10 9 21 21 nmos_a L=2.4e-07 W=1.2e-06 AD=7.2e-13 AS=4.8e-13 PD=1.8e-06 PS=9e-07 w_cont=6e-07 nfing=1 source_num=2 $X=51200 $Y=328060 $D=1
M7 9 12 gnd! gnd! nmos_a L=2.4e-07 W=1.2e-06 AD=7.2e-13 AS=4.8e-13 PD=1.8e-06 PS=9e-07 w_cont=6e-07 nfing=1 source_num=2 $X=56340 $Y=328040 $D=1
M8 12 nClk gnd! gnd! nmos_a L=2.4e-07 W=1.2e-06 AD=7.2e-13 AS=4.8e-13 PD=1.8e-06 PS=9e-07 w_cont=6e-07 nfing=1 source_num=2 $X=57780 $Y=328540 $D=1
M9 13 28 gnd! gnd! nmos_a L=2.4e-07 W=4.8e-07 AD=4.32e-13 AS=1.92e-13 PD=1.08e-06 PS=5.4e-07 w_cont=6e-07 nfing=1 source_num=2 $X=9180 $Y=329540 $D=1
M10 15 11 gnd! gnd! nmos_a L=2.4e-07 W=4.8e-07 AD=4.32e-13 AS=1.92e-13 PD=1.08e-06 PS=5.4e-07 w_cont=6e-07 nfing=1 source_num=2 $X=10600 $Y=327320 $D=1
M11 17 13 15 15 nmos_a L=2.4e-07 W=4.8e-07 AD=4.32e-13 AS=1.92e-13 PD=1.08e-06 PS=5.4e-07 w_cont=6e-07 nfing=1 source_num=2 $X=11300 $Y=329280 $D=1
M12 8 13 gnd! gnd! nmos_a L=2.4e-07 W=4.8e-07 AD=4.32e-13 AS=1.92e-13 PD=1.08e-06 PS=5.4e-07 w_cont=6e-07 nfing=1 source_num=2 $X=12040 $Y=327320 $D=1
M13 17 8 19 19 nmos_a L=2.4e-07 W=4.8e-07 AD=4.32e-13 AS=1.92e-13 PD=1.08e-06 PS=5.4e-07 w_cont=6e-07 nfing=1 source_num=2 $X=12700 $Y=329280 $D=1
M14 19 10 gnd! gnd! nmos_a L=2.4e-07 W=4.8e-07 AD=4.32e-13 AS=1.92e-13 PD=1.08e-06 PS=5.4e-07 w_cont=6e-07 nfing=1 source_num=2 $X=13520 $Y=327320 $D=1
M15 11 10 gnd! gnd! nmos_a L=2.4e-07 W=4.8e-07 AD=4.32e-13 AS=2.496e-13 PD=1.08e-06 PS=5.4e-07 w_cont=6e-07 nfing=1 source_num=2 $X=53320 $Y=327400 $D=1
M16 23 11 gnd! gnd! nmos_a L=2.4e-07 W=4.8e-07 AD=4.32e-13 AS=2.496e-13 PD=1.08e-06 PS=5.4e-07 w_cont=6e-07 nfing=1 source_num=2 $X=54080 $Y=327400 $D=1
M17 10 12 23 23 nmos_a L=2.4e-07 W=4.8e-07 AD=4.32e-13 AS=1.92e-13 PD=1.08e-06 PS=5.4e-07 w_cont=6e-07 nfing=1 source_num=2 $X=54940 $Y=328880 $D=1
M18 WEN 20 gnd! gnd! nmos_a L=2.4e-07 W=3.6e-06 AD=1.0816e-12 AS=1.44e-12 PD=2.08e-06 PS=2.08e-06 w_cont=1.6e-06 nfing=1 source_num=2 $X=28800 $Y=328040 $D=1
M19 WEN 20 gnd! gnd! nmos_a L=2.4e-07 W=3.6e-06 AD=1.0816e-12 AS=1.44e-12 PD=2.08e-06 PS=2.08e-06 w_cont=1.6e-06 nfing=1 source_num=2 $X=29560 $Y=328040 $D=1
M20 16 10 vdd! vdd! pmos_a L=2.4e-07 W=1e-06 AD=6.4e-13 AS=1.25e-13 PD=1.6e-06 PS=8e-07 w_cont=6e-07 nfing=1 mmm=1 $X=10540 $Y=333500 $D=5
M21 17 13 16 16 pmos_a L=2.4e-07 W=1e-06 AD=6.4e-13 AS=1.25e-13 PD=1.6e-06 PS=8e-07 w_cont=6e-07 nfing=1 mmm=1 $X=11300 $Y=331240 $D=5
M22 8 13 vdd! vdd! pmos_a L=2.4e-07 W=1e-06 AD=6.4e-13 AS=1.25e-13 PD=1.6e-06 PS=8e-07 w_cont=6e-07 nfing=1 mmm=1 $X=11980 $Y=333500 $D=5
M23 17 8 18 18 pmos_a L=2.4e-07 W=1e-06 AD=6.4e-13 AS=1.25e-13 PD=1.6e-06 PS=8e-07 w_cont=6e-07 nfing=1 mmm=1 $X=12700 $Y=331240 $D=5
M24 18 11 vdd! vdd! pmos_a L=2.4e-07 W=1e-06 AD=6.4e-13 AS=1.25e-13 PD=1.6e-06 PS=8e-07 w_cont=6e-07 nfing=1 mmm=1 $X=13420 $Y=333500 $D=5
M25 24 11 vdd! vdd! pmos_a L=2.4e-07 W=1e-06 AD=6.4e-13 AS=1.25e-13 PD=1.6e-06 PS=8e-07 w_cont=6e-07 nfing=1 mmm=1 $X=54080 $Y=333380 $D=5
M26 27 13 vdd! vdd! pmos_a L=2.4e-07 W=2e-06 AD=1.04e-12 AS=1.3e-13 PD=2.6e-06 PS=1.3e-06 w_cont=6e-07 nfing=1 mmm=1 $X=62300 $Y=331900 $D=5
M27 27 12 vdd! vdd! pmos_a L=2.4e-07 W=2e-06 AD=1.04e-12 AS=1.3e-13 PD=2.6e-06 PS=1.3e-06 w_cont=6e-07 nfing=1 mmm=1 $X=63740 $Y=331900 $D=5
M28 WEN 20 vdd! vdd! pmos_a L=2.4e-07 W=5.76e-06 AD=1.7836e-12 AS=2.488e-13 PD=3.43e-06 PS=3.43e-06 w_cont=1.1e-06 nfing=1 mmm=1 $X=31040 $Y=327380 $D=5
M29 WEN 20 vdd! vdd! pmos_a L=2.4e-07 W=5.76e-06 AD=1.7836e-12 AS=2.488e-13 PD=3.43e-06 PS=3.43e-06 w_cont=1.1e-06 nfing=1 mmm=1 $X=31800 $Y=327380 $D=5
M30 14 27 vdd! vdd! pmos_a L=2.4e-07 W=5.76e-06 AD=1.7836e-12 AS=2.488e-13 PD=3.43e-06 PS=3.43e-06 w_cont=1.1e-06 nfing=1 mmm=1 $X=67500 $Y=327340 $D=5
M31 14 27 vdd! vdd! pmos_a L=2.4e-07 W=5.76e-06 AD=1.7836e-12 AS=2.488e-13 PD=3.43e-06 PS=3.43e-06 w_cont=1.1e-06 nfing=1 mmm=1 $X=68260 $Y=327340 $D=5
M32 nWE 14 vdd! vdd! pmos_a L=2.4e-07 W=5.76e-06 AD=2.744e-12 AS=2.488e-13 PD=6.86e-06 PS=3.43e-06 w_cont=1.1e-06 nfing=1 mmm=1 $X=72940 $Y=327060 $D=5
M33 nWE 14 vdd! vdd! pmos_a L=2.4e-07 W=5.76e-06 AD=2.744e-12 AS=2.488e-13 PD=6.86e-06 PS=3.43e-06 w_cont=1.1e-06 nfing=1 mmm=1 $X=75780 $Y=327340 $D=5
M34 nWE 14 vdd! vdd! pmos_a L=2.4e-07 W=5.76e-06 AD=2.744e-12 AS=2.488e-13 PD=6.86e-06 PS=3.43e-06 w_cont=1.1e-06 nfing=1 mmm=1 $X=80460 $Y=327060 $D=5
M35 nWE 14 vdd! vdd! pmos_a L=2.4e-07 W=5.76e-06 AD=2.744e-12 AS=2.488e-13 PD=6.86e-06 PS=3.43e-06 w_cont=1.1e-06 nfing=1 mmm=1 $X=83300 $Y=327340 $D=5
M36 nWE 14 vdd! vdd! pmos_a L=2.4e-07 W=5.76e-06 AD=2.744e-12 AS=2.488e-13 PD=6.86e-06 PS=3.43e-06 w_cont=1.1e-06 nfing=1 mmm=1 $X=87980 $Y=327060 $D=5
M37 nWE 14 vdd! vdd! pmos_a L=2.4e-07 W=5.76e-06 AD=2.744e-12 AS=2.488e-13 PD=6.86e-06 PS=3.43e-06 w_cont=1.1e-06 nfing=1 mmm=1 $X=90820 $Y=327340 $D=5
M38 nWE 14 vdd! vdd! pmos_a L=2.4e-07 W=5.76e-06 AD=2.744e-12 AS=2.488e-13 PD=6.86e-06 PS=3.43e-06 w_cont=1.1e-06 nfing=1 mmm=1 $X=95500 $Y=327060 $D=5
M39 nWE 14 vdd! vdd! pmos_a L=2.4e-07 W=5.76e-06 AD=2.744e-12 AS=2.488e-13 PD=6.86e-06 PS=3.43e-06 w_cont=1.1e-06 nfing=1 mmm=1 $X=98340 $Y=327340 $D=5
M40 nATD 17 vdd! vdd! pmos_a L=2.4e-07 W=2e-06 AD=1.04e-12 AS=1.3e-13 PD=2.6e-06 PS=1.3e-06 w_cont=6e-07 nfing=1 mmm=1 $X=14960 $Y=331120 $D=5
M41 20 8 vdd! vdd! pmos_a L=2.4e-07 W=2e-06 AD=1.04e-12 AS=1.3e-13 PD=2.6e-06 PS=1.3e-06 w_cont=6e-07 nfing=1 mmm=1 $X=27360 $Y=331300 $D=5
M42 22 13 vdd! vdd! pmos_a L=2.4e-07 W=2e-06 AD=1.04e-12 AS=1.3e-13 PD=2.6e-06 PS=1.3e-06 w_cont=6e-07 nfing=1 mmm=1 $X=49760 $Y=331200 $D=5
M43 10 12 22 22 pmos_a L=2.4e-07 W=2e-06 AD=1.04e-12 AS=1.3e-13 PD=2.6e-06 PS=1.3e-06 w_cont=6e-07 nfing=1 mmm=1 $X=51200 $Y=330880 $D=5
M44 9 12 vdd! vdd! pmos_a L=2.4e-07 W=2e-06 AD=1.04e-12 AS=1.3e-13 PD=2.6e-06 PS=1.3e-06 w_cont=6e-07 nfing=1 mmm=1 $X=56340 $Y=330240 $D=5
M45 12 nClk vdd! vdd! pmos_a L=2.4e-07 W=2e-06 AD=1.04e-12 AS=1.3e-13 PD=2.6e-06 PS=1.3e-06 w_cont=6e-07 nfing=1 mmm=1 $X=57780 $Y=331820 $D=5
M46 27 11 vdd! vdd! pmos_a L=2.4e-07 W=2e-06 AD=1.04e-12 AS=1.3e-13 PD=2.6e-06 PS=1.3e-06 w_cont=6e-07 nfing=1 mmm=1 $X=60860 $Y=331900 $D=5
M47 11 10 vdd! vdd! pmos_a L=2.4e-07 W=1e-06 AD=6.4e-13 AS=1.25e-13 PD=1.6e-06 PS=8e-07 w_cont=6e-07 nfing=1 mmm=1 $X=52640 $Y=332380 $D=5
M48 10 9 24 24 pmos_a L=2.4e-07 W=1e-06 AD=6.4e-13 AS=1.25e-13 PD=1.6e-06 PS=8e-07 w_cont=6e-07 nfing=1 mmm=1 $X=54940 $Y=331320 $D=5
M49 13 28 vdd! vdd! pmos_a L=2.4e-07 W=4.8e-07 AD=4.32e-13 AS=1.224e-13 PD=1.08e-06 PS=5.4e-07 w_cont=6e-07 nfing=1 mmm=1 $X=9180 $Y=331600 $D=5
M50 vdd! gnd! vdd! cpoly_n w=6e-06 l=2e-06 c=7.5402e-14 as=2.4e-13 ad=2.304e-12 ps=2.88e-06 pd=4.86761e-06 sim_w=5.76e-06 m_per_maxw=1.04167 numb_sub_cont=3 nfing=1 $X=36160 $Y=328200 $D=22
M51 vdd! gnd! vdd! cpoly_n w=6e-06 l=2e-06 c=7.5402e-14 as=2.4e-13 ad=2.304e-12 ps=2.88e-06 pd=4.86761e-06 sim_w=5.76e-06 m_per_maxw=1.04167 numb_sub_cont=3 nfing=1 $X=43680 $Y=328200 $D=22
M52 vdd! gnd! vdd! cpoly_n w=6e-06 l=2e-06 c=7.5402e-14 as=2.4e-13 ad=2.304e-12 ps=2.88e-06 pd=4.86761e-06 sim_w=5.76e-06 m_per_maxw=1.04167 numb_sub_cont=3 nfing=1 $X=69740 $Y=328200 $D=22
M53 vdd! gnd! vdd! cpoly_n w=6e-06 l=2e-06 c=7.5402e-14 as=2.4e-13 ad=2.304e-12 ps=2.88e-06 pd=4.86761e-06 sim_w=5.76e-06 m_per_maxw=1.04167 numb_sub_cont=3 nfing=1 $X=77260 $Y=328200 $D=22
M54 vdd! gnd! vdd! cpoly_n w=6e-06 l=2e-06 c=7.5402e-14 as=2.4e-13 ad=2.304e-12 ps=2.88e-06 pd=4.86761e-06 sim_w=5.76e-06 m_per_maxw=1.04167 numb_sub_cont=3 nfing=1 $X=84780 $Y=328200 $D=22
M55 vdd! gnd! vdd! cpoly_n w=6e-06 l=2e-06 c=7.5402e-14 as=2.4e-13 ad=2.304e-12 ps=2.88e-06 pd=4.86761e-06 sim_w=5.76e-06 m_per_maxw=1.04167 numb_sub_cont=3 nfing=1 $X=92300 $Y=328200 $D=22
D56 NWR vdd! dn PJ=0.0002 m=1 $X=4020 $Y=-95300 $D=9
D57 NWR vdd! dn PJ=0.0002 m=1 $X=4020 $Y=114700 $D=9
D58 gnd! NWR dn PJ=0.0002 m=1 $X=6340 $Y=-99700 $D=9
D59 gnd! NWR dn PJ=0.0002 m=1 $X=6340 $Y=110300 $D=9
D60 NWR vdd! dn PJ=0.0002 m=1 $X=8660 $Y=-95300 $D=9
D61 NWR vdd! dn PJ=0.0002 m=1 $X=8660 $Y=114700 $D=9
D62 gnd! NWR dn PJ=0.0001 m=1 $X=10980 $Y=-99700 $D=9
D63 gnd! NWR dn PJ=0.0001 m=1 $X=10980 $Y=110300 $D=9
D64 NWR vdd! dn PJ=0.0001 m=1 $X=14160 $Y=4700 $D=9
D65 NWR vdd! dn PJ=0.0001 m=1 $X=14160 $Y=214700 $D=9
D66 gnd! NWR dn PJ=0.0002 m=1 $X=16480 $Y=-99700 $D=9
D67 gnd! NWR dn PJ=0.0002 m=1 $X=16480 $Y=110300 $D=9
D68 NWR vdd! dn PJ=0.0002 m=1 $X=18800 $Y=-95300 $D=9
D69 NWR vdd! dn PJ=0.0002 m=1 $X=18800 $Y=114700 $D=9
D70 gnd! NWR dn PJ=0.0002 m=1 $X=21120 $Y=-99700 $D=9
D71 gnd! NWR dn PJ=0.0002 m=1 $X=21120 $Y=110300 $D=9
D72 NWR vdd! dn PJ=0.0002 m=1 $X=23440 $Y=-95300 $D=9
D73 NWR vdd! dn PJ=0.0002 m=1 $X=23440 $Y=114700 $D=9
D74 gnd! NWR dn PJ=0.0001 m=1 $X=25760 $Y=-99700 $D=9
D75 gnd! NWR dn PJ=0.0001 m=1 $X=25760 $Y=110300 $D=9
D76 NWR vdd! dn PJ=0.0001 m=1 $X=28940 $Y=4700 $D=9
D77 NWR vdd! dn PJ=0.0001 m=1 $X=28940 $Y=214700 $D=9
D78 gnd! NWR dn PJ=0.0002 m=1 $X=31260 $Y=-99700 $D=9
D79 gnd! NWR dn PJ=0.0002 m=1 $X=31260 $Y=110300 $D=9
D80 NWR vdd! dn PJ=0.0002 m=1 $X=33580 $Y=-95300 $D=9
D81 NWR vdd! dn PJ=0.0002 m=1 $X=33580 $Y=114700 $D=9
D82 gnd! NWR dn PJ=0.0002 m=1 $X=35900 $Y=-99700 $D=9
D83 gnd! NWR dn PJ=0.0002 m=1 $X=35900 $Y=110300 $D=9
D84 NWR vdd! dn PJ=0.0002 m=1 $X=38220 $Y=-95300 $D=9
D85 NWR vdd! dn PJ=0.0002 m=1 $X=38220 $Y=114700 $D=9
D86 gnd! NWR dn PJ=0.0001 m=1 $X=40540 $Y=-99700 $D=9
D87 gnd! NWR dn PJ=0.0001 m=1 $X=40540 $Y=110300 $D=9
D88 NWR vdd! dn PJ=0.0001 m=1 $X=43720 $Y=4700 $D=9
D89 NWR vdd! dn PJ=0.0001 m=1 $X=43720 $Y=214700 $D=9
D90 gnd! NWR dn PJ=0.0002 m=1 $X=46040 $Y=-99700 $D=9
D91 gnd! NWR dn PJ=0.0002 m=1 $X=46040 $Y=110300 $D=9
D92 NWR vdd! dn PJ=0.0002 m=1 $X=48360 $Y=-95300 $D=9
D93 NWR vdd! dn PJ=0.0002 m=1 $X=48360 $Y=114700 $D=9
D94 gnd! NWR dn PJ=0.0002 m=1 $X=50680 $Y=-99700 $D=9
D95 gnd! NWR dn PJ=0.0002 m=1 $X=50680 $Y=110300 $D=9
D96 NWR vdd! dn PJ=0.0002 m=1 $X=53000 $Y=-95300 $D=9
D97 NWR vdd! dn PJ=0.0002 m=1 $X=53000 $Y=114700 $D=9
D98 gnd! NWR dn PJ=0.0001 m=1 $X=55320 $Y=-99700 $D=9
D99 gnd! NWR dn PJ=0.0001 m=1 $X=55320 $Y=110300 $D=9
D100 NWR vdd! dn PJ=0.0001 m=1 $X=58500 $Y=4700 $D=9
D101 NWR vdd! dn PJ=0.0001 m=1 $X=58500 $Y=214700 $D=9
D102 gnd! NWR dn PJ=0.0002 m=1 $X=60820 $Y=-99700 $D=9
D103 gnd! NWR dn PJ=0.0002 m=1 $X=60820 $Y=110300 $D=9
D104 NWR vdd! dn PJ=0.0002 m=1 $X=63140 $Y=-95300 $D=9
D105 NWR vdd! dn PJ=0.0002 m=1 $X=63140 $Y=114700 $D=9
D106 gnd! NWR dn PJ=0.0002 m=1 $X=65460 $Y=-99700 $D=9
D107 gnd! NWR dn PJ=0.0002 m=1 $X=65460 $Y=110300 $D=9
D108 NWR vdd! dn PJ=0.0002 m=1 $X=67780 $Y=-95300 $D=9
D109 NWR vdd! dn PJ=0.0002 m=1 $X=67780 $Y=114700 $D=9
D110 gnd! NWR dn PJ=0.0001 m=1 $X=70100 $Y=-99700 $D=9
D111 gnd! NWR dn PJ=0.0001 m=1 $X=70100 $Y=110300 $D=9
D112 NWR vdd! dn PJ=0.0001 m=1 $X=73280 $Y=4700 $D=9
D113 NWR vdd! dn PJ=0.0001 m=1 $X=73280 $Y=214700 $D=9
D114 gnd! NWR dn PJ=0.0002 m=1 $X=75600 $Y=-99700 $D=9
D115 gnd! NWR dn PJ=0.0002 m=1 $X=75600 $Y=110300 $D=9
D116 NWR vdd! dn PJ=0.0002 m=1 $X=77920 $Y=-95300 $D=9
D117 NWR vdd! dn PJ=0.0002 m=1 $X=77920 $Y=114700 $D=9
D118 gnd! NWR dn PJ=0.0002 m=1 $X=80240 $Y=-99700 $D=9
D119 gnd! NWR dn PJ=0.0002 m=1 $X=80240 $Y=110300 $D=9
D120 NWR vdd! dn PJ=0.0002 m=1 $X=82560 $Y=-95300 $D=9
D121 NWR vdd! dn PJ=0.0002 m=1 $X=82560 $Y=114700 $D=9
D122 gnd! NWR dn PJ=0.0001 m=1 $X=84880 $Y=-99700 $D=9
D123 gnd! NWR dn PJ=0.0001 m=1 $X=84880 $Y=110300 $D=9
D124 NWR vdd! dn PJ=0.0001 m=1 $X=88060 $Y=4700 $D=9
D125 NWR vdd! dn PJ=0.0001 m=1 $X=88060 $Y=214700 $D=9
D126 gnd! NWR dn PJ=0.0002 m=1 $X=90380 $Y=-99700 $D=9
D127 gnd! NWR dn PJ=0.0002 m=1 $X=90380 $Y=110300 $D=9
D128 NWR vdd! dn PJ=0.0002 m=1 $X=92700 $Y=-95300 $D=9
D129 NWR vdd! dn PJ=0.0002 m=1 $X=92700 $Y=114700 $D=9
D130 gnd! NWR dn PJ=0.0002 m=1 $X=95020 $Y=-99700 $D=9
D131 gnd! NWR dn PJ=0.0002 m=1 $X=95020 $Y=110300 $D=9
D132 gnd! 28 dn PJ=5e-06 m=1 $X=1560 $Y=328560 $D=10
D133 28 vdd! dn PJ=5e-06 m=1 $X=1560 $Y=334960 $D=10
D134 gnd! 28 dn PJ=5e-06 m=1 $X=1560 $Y=329900 $D=11
D135 28 vdd! dn PJ=5e-06 m=1 $X=1560 $Y=332220 $D=11
X151 gnd! 14 27 nmos_a_CDNS_5887047866553 $T=65440 327140 0 0 $X=65440 $Y=327140
X152 gnd! nWE 14 nmos_a_CDNS_5887047866553 $T=73760 327140 0 0 $X=73760 $Y=327140
X153 gnd! nWE 14 nmos_a_CDNS_5887047866553 $T=81280 327140 0 0 $X=81280 $Y=327140
X154 gnd! nWE 14 nmos_a_CDNS_5887047866553 $T=88800 327140 0 0 $X=88800 $Y=327140
X155 gnd! nWE 14 nmos_a_CDNS_5887047866553 $T=96320 327140 0 0 $X=96320 $Y=327140
X189 gnd! vdd! cpoly_p_CDNS_5887047866511 $T=7980 317780 0 0 $X=7980 $Y=317780
X190 vdd! gnd! cpoly_n_CDNS_5887047866514 $T=520 336500 0 0 $X=520 $Y=336500
X191 NWR 28 PAD $T=0 1440 0 0 $X=-5000 $Y=-235000
.ENDS
***************************************
.SUBCKT cpoly_p_CDNS_58870478665105 1 2
** N=2 EP=2 IP=0 FDC=62
M0 1 2 1 cpoly_p w=8.62e-06 l=2e-06 c=1.08536e-13 as=1.21314e-13 ad=7.488e-13 ps=1.44e-06 pd=1.21456e-06 sim_w=2.88e-06 m_per_maxw=2.99306 numb_sub_cont=4 nfing=1 $X=620 $Y=200 $D=21
M1 1 2 1 cpoly_p w=8.62e-06 l=2e-06 c=1.08536e-13 as=1.53388e-13 ad=7.488e-13 ps=1.44e-06 pd=1.21456e-06 sim_w=2.88e-06 m_per_maxw=2.99306 numb_sub_cont=4 nfing=1 $X=3140 $Y=200 $D=21
M2 1 2 1 cpoly_p w=8.62e-06 l=2e-06 c=1.08536e-13 as=1.53388e-13 ad=7.488e-13 ps=1.44e-06 pd=1.21456e-06 sim_w=2.88e-06 m_per_maxw=2.99306 numb_sub_cont=4 nfing=1 $X=5660 $Y=200 $D=21
M3 1 2 1 cpoly_p w=8.62e-06 l=2e-06 c=1.08536e-13 as=1.53388e-13 ad=7.488e-13 ps=1.44e-06 pd=1.21456e-06 sim_w=2.88e-06 m_per_maxw=2.99306 numb_sub_cont=4 nfing=1 $X=8180 $Y=200 $D=21
M4 1 2 1 cpoly_p w=8.62e-06 l=2e-06 c=1.08536e-13 as=1.53388e-13 ad=7.488e-13 ps=1.44e-06 pd=1.21456e-06 sim_w=2.88e-06 m_per_maxw=2.99306 numb_sub_cont=4 nfing=1 $X=10700 $Y=200 $D=21
M5 1 2 1 cpoly_p w=8.62e-06 l=2e-06 c=1.08536e-13 as=1.53388e-13 ad=7.488e-13 ps=1.44e-06 pd=1.21456e-06 sim_w=2.88e-06 m_per_maxw=2.99306 numb_sub_cont=4 nfing=1 $X=13220 $Y=200 $D=21
M6 1 2 1 cpoly_p w=8.62e-06 l=2e-06 c=1.08536e-13 as=1.53388e-13 ad=7.488e-13 ps=1.44e-06 pd=1.21456e-06 sim_w=2.88e-06 m_per_maxw=2.99306 numb_sub_cont=4 nfing=1 $X=15740 $Y=200 $D=21
M7 1 2 1 cpoly_p w=8.62e-06 l=2e-06 c=1.08536e-13 as=1.53388e-13 ad=7.488e-13 ps=1.44e-06 pd=1.21456e-06 sim_w=2.88e-06 m_per_maxw=2.99306 numb_sub_cont=4 nfing=1 $X=18260 $Y=200 $D=21
M8 1 2 1 cpoly_p w=8.62e-06 l=2e-06 c=1.08536e-13 as=1.53388e-13 ad=7.488e-13 ps=1.44e-06 pd=1.21456e-06 sim_w=2.88e-06 m_per_maxw=2.99306 numb_sub_cont=4 nfing=1 $X=20780 $Y=200 $D=21
M9 1 2 1 cpoly_p w=8.62e-06 l=2e-06 c=1.08536e-13 as=1.53388e-13 ad=7.488e-13 ps=1.44e-06 pd=1.21456e-06 sim_w=2.88e-06 m_per_maxw=2.99306 numb_sub_cont=4 nfing=1 $X=23300 $Y=200 $D=21
M10 1 2 1 cpoly_p w=8.62e-06 l=2e-06 c=1.08536e-13 as=1.53388e-13 ad=7.488e-13 ps=1.44e-06 pd=1.21456e-06 sim_w=2.88e-06 m_per_maxw=2.99306 numb_sub_cont=4 nfing=1 $X=25820 $Y=200 $D=21
M11 1 2 1 cpoly_p w=8.62e-06 l=2e-06 c=1.08536e-13 as=1.53388e-13 ad=7.488e-13 ps=1.44e-06 pd=1.21456e-06 sim_w=2.88e-06 m_per_maxw=2.99306 numb_sub_cont=4 nfing=1 $X=28340 $Y=200 $D=21
M12 1 2 1 cpoly_p w=8.62e-06 l=2e-06 c=1.08536e-13 as=1.53388e-13 ad=7.488e-13 ps=1.44e-06 pd=1.21456e-06 sim_w=2.88e-06 m_per_maxw=2.99306 numb_sub_cont=4 nfing=1 $X=30860 $Y=200 $D=21
M13 1 2 1 cpoly_p w=8.62e-06 l=2e-06 c=1.08536e-13 as=1.53388e-13 ad=7.488e-13 ps=1.44e-06 pd=1.21456e-06 sim_w=2.88e-06 m_per_maxw=2.99306 numb_sub_cont=4 nfing=1 $X=33380 $Y=200 $D=21
M14 1 2 1 cpoly_p w=8.62e-06 l=2e-06 c=1.08536e-13 as=1.53388e-13 ad=7.488e-13 ps=1.44e-06 pd=1.21456e-06 sim_w=2.88e-06 m_per_maxw=2.99306 numb_sub_cont=4 nfing=1 $X=35900 $Y=200 $D=21
M15 1 2 1 cpoly_p w=8.62e-06 l=2e-06 c=1.08536e-13 as=1.53388e-13 ad=7.488e-13 ps=1.44e-06 pd=1.21456e-06 sim_w=2.88e-06 m_per_maxw=2.99306 numb_sub_cont=4 nfing=1 $X=38420 $Y=200 $D=21
M16 1 2 1 cpoly_p w=8.62e-06 l=2e-06 c=1.08536e-13 as=1.53388e-13 ad=7.488e-13 ps=1.44e-06 pd=1.21456e-06 sim_w=2.88e-06 m_per_maxw=2.99306 numb_sub_cont=4 nfing=1 $X=40940 $Y=200 $D=21
M17 1 2 1 cpoly_p w=8.62e-06 l=2e-06 c=1.08536e-13 as=1.53388e-13 ad=7.488e-13 ps=1.44e-06 pd=1.21456e-06 sim_w=2.88e-06 m_per_maxw=2.99306 numb_sub_cont=4 nfing=1 $X=43460 $Y=200 $D=21
M18 1 2 1 cpoly_p w=8.62e-06 l=2e-06 c=1.08536e-13 as=1.53388e-13 ad=7.488e-13 ps=1.44e-06 pd=1.21456e-06 sim_w=2.88e-06 m_per_maxw=2.99306 numb_sub_cont=4 nfing=1 $X=45980 $Y=200 $D=21
M19 1 2 1 cpoly_p w=8.62e-06 l=2e-06 c=1.08536e-13 as=1.53388e-13 ad=7.488e-13 ps=1.44e-06 pd=1.21456e-06 sim_w=2.88e-06 m_per_maxw=2.99306 numb_sub_cont=4 nfing=1 $X=48500 $Y=200 $D=21
M20 1 2 1 cpoly_p w=8.62e-06 l=2e-06 c=1.08536e-13 as=1.53388e-13 ad=7.488e-13 ps=1.44e-06 pd=1.21456e-06 sim_w=2.88e-06 m_per_maxw=2.99306 numb_sub_cont=4 nfing=1 $X=51020 $Y=200 $D=21
M21 1 2 1 cpoly_p w=8.62e-06 l=2e-06 c=1.08536e-13 as=1.53388e-13 ad=7.488e-13 ps=1.44e-06 pd=1.21456e-06 sim_w=2.88e-06 m_per_maxw=2.99306 numb_sub_cont=4 nfing=1 $X=53540 $Y=200 $D=21
M22 1 2 1 cpoly_p w=8.62e-06 l=2e-06 c=1.08536e-13 as=1.53388e-13 ad=7.488e-13 ps=1.44e-06 pd=1.21456e-06 sim_w=2.88e-06 m_per_maxw=2.99306 numb_sub_cont=4 nfing=1 $X=56060 $Y=200 $D=21
M23 1 2 1 cpoly_p w=8.62e-06 l=2e-06 c=1.08536e-13 as=1.53388e-13 ad=7.488e-13 ps=1.44e-06 pd=1.21456e-06 sim_w=2.88e-06 m_per_maxw=2.99306 numb_sub_cont=4 nfing=1 $X=58580 $Y=200 $D=21
M24 1 2 1 cpoly_p w=8.62e-06 l=2e-06 c=1.08536e-13 as=1.53388e-13 ad=7.488e-13 ps=1.44e-06 pd=1.21456e-06 sim_w=2.88e-06 m_per_maxw=2.99306 numb_sub_cont=4 nfing=1 $X=61100 $Y=200 $D=21
M25 1 2 1 cpoly_p w=8.62e-06 l=2e-06 c=1.08536e-13 as=1.53388e-13 ad=7.488e-13 ps=1.44e-06 pd=1.21456e-06 sim_w=2.88e-06 m_per_maxw=2.99306 numb_sub_cont=4 nfing=1 $X=63620 $Y=200 $D=21
M26 1 2 1 cpoly_p w=8.62e-06 l=2e-06 c=1.08536e-13 as=1.53388e-13 ad=7.488e-13 ps=1.44e-06 pd=1.21456e-06 sim_w=2.88e-06 m_per_maxw=2.99306 numb_sub_cont=4 nfing=1 $X=66140 $Y=200 $D=21
M27 1 2 1 cpoly_p w=8.62e-06 l=2e-06 c=1.08536e-13 as=1.53388e-13 ad=7.488e-13 ps=1.44e-06 pd=1.21456e-06 sim_w=2.88e-06 m_per_maxw=2.99306 numb_sub_cont=4 nfing=1 $X=68660 $Y=200 $D=21
M28 1 2 1 cpoly_p w=8.62e-06 l=2e-06 c=1.08536e-13 as=1.53388e-13 ad=7.488e-13 ps=1.44e-06 pd=1.21456e-06 sim_w=2.88e-06 m_per_maxw=2.99306 numb_sub_cont=4 nfing=1 $X=71180 $Y=200 $D=21
M29 1 2 1 cpoly_p w=8.62e-06 l=2e-06 c=1.08536e-13 as=1.53388e-13 ad=7.488e-13 ps=1.44e-06 pd=1.21456e-06 sim_w=2.88e-06 m_per_maxw=2.99306 numb_sub_cont=4 nfing=1 $X=73700 $Y=200 $D=21
M30 1 2 1 cpoly_p w=8.62e-06 l=2e-06 c=1.08536e-13 as=1.53388e-13 ad=7.488e-13 ps=1.44e-06 pd=1.21456e-06 sim_w=2.88e-06 m_per_maxw=2.99306 numb_sub_cont=4 nfing=1 $X=76220 $Y=200 $D=21
M31 1 2 1 cpoly_p w=8.62e-06 l=2e-06 c=1.08536e-13 as=1.53388e-13 ad=7.488e-13 ps=1.44e-06 pd=1.21456e-06 sim_w=2.88e-06 m_per_maxw=2.99306 numb_sub_cont=4 nfing=1 $X=78740 $Y=200 $D=21
M32 1 2 1 cpoly_p w=8.62e-06 l=2e-06 c=1.08536e-13 as=1.53388e-13 ad=7.488e-13 ps=1.44e-06 pd=1.21456e-06 sim_w=2.88e-06 m_per_maxw=2.99306 numb_sub_cont=4 nfing=1 $X=81260 $Y=200 $D=21
M33 1 2 1 cpoly_p w=8.62e-06 l=2e-06 c=1.08536e-13 as=1.53388e-13 ad=7.488e-13 ps=1.44e-06 pd=1.21456e-06 sim_w=2.88e-06 m_per_maxw=2.99306 numb_sub_cont=4 nfing=1 $X=83780 $Y=200 $D=21
M34 1 2 1 cpoly_p w=8.62e-06 l=2e-06 c=1.08536e-13 as=1.53388e-13 ad=7.488e-13 ps=1.44e-06 pd=1.21456e-06 sim_w=2.88e-06 m_per_maxw=2.99306 numb_sub_cont=4 nfing=1 $X=86300 $Y=200 $D=21
M35 1 2 1 cpoly_p w=8.62e-06 l=2e-06 c=1.08536e-13 as=1.53388e-13 ad=7.488e-13 ps=1.44e-06 pd=1.21456e-06 sim_w=2.88e-06 m_per_maxw=2.99306 numb_sub_cont=4 nfing=1 $X=88820 $Y=200 $D=21
M36 1 2 1 cpoly_p w=8.62e-06 l=2e-06 c=1.08536e-13 as=1.53388e-13 ad=7.488e-13 ps=1.44e-06 pd=1.21456e-06 sim_w=2.88e-06 m_per_maxw=2.99306 numb_sub_cont=4 nfing=1 $X=91340 $Y=200 $D=21
M37 1 2 1 cpoly_p w=8.62e-06 l=2e-06 c=1.08536e-13 as=1.53388e-13 ad=7.488e-13 ps=1.44e-06 pd=1.21456e-06 sim_w=2.88e-06 m_per_maxw=2.99306 numb_sub_cont=4 nfing=1 $X=93860 $Y=200 $D=21
M38 1 2 1 cpoly_p w=8.62e-06 l=2e-06 c=1.08536e-13 as=1.53388e-13 ad=7.488e-13 ps=1.44e-06 pd=1.21456e-06 sim_w=2.88e-06 m_per_maxw=2.99306 numb_sub_cont=4 nfing=1 $X=96380 $Y=200 $D=21
M39 1 2 1 cpoly_p w=8.62e-06 l=2e-06 c=1.08536e-13 as=1.53388e-13 ad=7.488e-13 ps=1.44e-06 pd=1.21456e-06 sim_w=2.88e-06 m_per_maxw=2.99306 numb_sub_cont=4 nfing=1 $X=98900 $Y=200 $D=21
M40 1 2 1 cpoly_p w=8.62e-06 l=2e-06 c=1.08536e-13 as=1.53388e-13 ad=7.488e-13 ps=1.44e-06 pd=1.21456e-06 sim_w=2.88e-06 m_per_maxw=2.99306 numb_sub_cont=4 nfing=1 $X=101420 $Y=200 $D=21
M41 1 2 1 cpoly_p w=8.62e-06 l=2e-06 c=1.08536e-13 as=1.53388e-13 ad=7.488e-13 ps=1.44e-06 pd=1.21456e-06 sim_w=2.88e-06 m_per_maxw=2.99306 numb_sub_cont=4 nfing=1 $X=103940 $Y=200 $D=21
M42 1 2 1 cpoly_p w=8.62e-06 l=2e-06 c=1.08536e-13 as=1.53388e-13 ad=7.488e-13 ps=1.44e-06 pd=1.21456e-06 sim_w=2.88e-06 m_per_maxw=2.99306 numb_sub_cont=4 nfing=1 $X=106460 $Y=200 $D=21
M43 1 2 1 cpoly_p w=8.62e-06 l=2e-06 c=1.08536e-13 as=1.53388e-13 ad=7.488e-13 ps=1.44e-06 pd=1.21456e-06 sim_w=2.88e-06 m_per_maxw=2.99306 numb_sub_cont=4 nfing=1 $X=108980 $Y=200 $D=21
M44 1 2 1 cpoly_p w=8.62e-06 l=2e-06 c=1.08536e-13 as=1.53388e-13 ad=7.488e-13 ps=1.44e-06 pd=1.21456e-06 sim_w=2.88e-06 m_per_maxw=2.99306 numb_sub_cont=4 nfing=1 $X=111500 $Y=200 $D=21
M45 1 2 1 cpoly_p w=8.62e-06 l=2e-06 c=1.08536e-13 as=1.53388e-13 ad=7.488e-13 ps=1.44e-06 pd=1.21456e-06 sim_w=2.88e-06 m_per_maxw=2.99306 numb_sub_cont=4 nfing=1 $X=114020 $Y=200 $D=21
M46 1 2 1 cpoly_p w=8.62e-06 l=2e-06 c=1.08536e-13 as=1.53388e-13 ad=7.488e-13 ps=1.44e-06 pd=1.21456e-06 sim_w=2.88e-06 m_per_maxw=2.99306 numb_sub_cont=4 nfing=1 $X=116540 $Y=200 $D=21
M47 1 2 1 cpoly_p w=8.62e-06 l=2e-06 c=1.08536e-13 as=1.53388e-13 ad=7.488e-13 ps=1.44e-06 pd=1.21456e-06 sim_w=2.88e-06 m_per_maxw=2.99306 numb_sub_cont=4 nfing=1 $X=119060 $Y=200 $D=21
M48 1 2 1 cpoly_p w=8.62e-06 l=2e-06 c=1.08536e-13 as=1.53388e-13 ad=7.488e-13 ps=1.44e-06 pd=1.21456e-06 sim_w=2.88e-06 m_per_maxw=2.99306 numb_sub_cont=4 nfing=1 $X=121580 $Y=200 $D=21
M49 1 2 1 cpoly_p w=8.62e-06 l=2e-06 c=1.08536e-13 as=1.53388e-13 ad=7.488e-13 ps=1.44e-06 pd=1.21456e-06 sim_w=2.88e-06 m_per_maxw=2.99306 numb_sub_cont=4 nfing=1 $X=124100 $Y=200 $D=21
M50 1 2 1 cpoly_p w=8.62e-06 l=2e-06 c=1.08536e-13 as=1.53388e-13 ad=7.488e-13 ps=1.44e-06 pd=1.21456e-06 sim_w=2.88e-06 m_per_maxw=2.99306 numb_sub_cont=4 nfing=1 $X=126620 $Y=200 $D=21
M51 1 2 1 cpoly_p w=8.62e-06 l=2e-06 c=1.08536e-13 as=1.53388e-13 ad=7.488e-13 ps=1.44e-06 pd=1.21456e-06 sim_w=2.88e-06 m_per_maxw=2.99306 numb_sub_cont=4 nfing=1 $X=129140 $Y=200 $D=21
M52 1 2 1 cpoly_p w=8.62e-06 l=2e-06 c=1.08536e-13 as=1.53388e-13 ad=7.488e-13 ps=1.44e-06 pd=1.21456e-06 sim_w=2.88e-06 m_per_maxw=2.99306 numb_sub_cont=4 nfing=1 $X=131660 $Y=200 $D=21
M53 1 2 1 cpoly_p w=8.62e-06 l=2e-06 c=1.08536e-13 as=1.53388e-13 ad=7.488e-13 ps=1.44e-06 pd=1.21456e-06 sim_w=2.88e-06 m_per_maxw=2.99306 numb_sub_cont=4 nfing=1 $X=134180 $Y=200 $D=21
M54 1 2 1 cpoly_p w=8.62e-06 l=2e-06 c=1.08536e-13 as=1.53388e-13 ad=7.488e-13 ps=1.44e-06 pd=1.21456e-06 sim_w=2.88e-06 m_per_maxw=2.99306 numb_sub_cont=4 nfing=1 $X=136700 $Y=200 $D=21
M55 1 2 1 cpoly_p w=8.62e-06 l=2e-06 c=1.08536e-13 as=1.53388e-13 ad=7.488e-13 ps=1.44e-06 pd=1.21456e-06 sim_w=2.88e-06 m_per_maxw=2.99306 numb_sub_cont=4 nfing=1 $X=139220 $Y=200 $D=21
M56 1 2 1 cpoly_p w=8.62e-06 l=2e-06 c=1.08536e-13 as=1.53388e-13 ad=7.488e-13 ps=1.44e-06 pd=1.21456e-06 sim_w=2.88e-06 m_per_maxw=2.99306 numb_sub_cont=4 nfing=1 $X=141740 $Y=200 $D=21
M57 1 2 1 cpoly_p w=8.62e-06 l=2e-06 c=1.08536e-13 as=1.53388e-13 ad=7.488e-13 ps=1.44e-06 pd=1.21456e-06 sim_w=2.88e-06 m_per_maxw=2.99306 numb_sub_cont=4 nfing=1 $X=144260 $Y=200 $D=21
M58 1 2 1 cpoly_p w=8.62e-06 l=2e-06 c=1.08536e-13 as=1.53388e-13 ad=7.488e-13 ps=1.44e-06 pd=1.21456e-06 sim_w=2.88e-06 m_per_maxw=2.99306 numb_sub_cont=4 nfing=1 $X=146780 $Y=200 $D=21
M59 1 2 1 cpoly_p w=8.62e-06 l=2e-06 c=1.08536e-13 as=1.53388e-13 ad=7.488e-13 ps=1.44e-06 pd=1.21456e-06 sim_w=2.88e-06 m_per_maxw=2.99306 numb_sub_cont=4 nfing=1 $X=149300 $Y=200 $D=21
M60 1 2 1 cpoly_p w=8.62e-06 l=2e-06 c=1.08536e-13 as=1.53388e-13 ad=7.488e-13 ps=1.44e-06 pd=1.21456e-06 sim_w=2.88e-06 m_per_maxw=2.99306 numb_sub_cont=4 nfing=1 $X=151820 $Y=200 $D=21
M61 1 2 1 cpoly_p w=8.62e-06 l=2e-06 c=1.08536e-13 as=1.21314e-13 ad=7.488e-13 ps=1.44e-06 pd=1.21456e-06 sim_w=2.88e-06 m_per_maxw=2.99306 numb_sub_cont=4 nfing=1 $X=154340 $Y=200 $D=21
.ENDS
***************************************
.SUBCKT cpoly_n_CDNS_58870478665104 1 2
** N=2 EP=2 IP=0 FDC=62
M0 1 2 1 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=1.67141e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=620 $Y=200 $D=22
M1 1 2 1 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=3140 $Y=200 $D=22
M2 1 2 1 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=5660 $Y=200 $D=22
M3 1 2 1 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=8180 $Y=200 $D=22
M4 1 2 1 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=10700 $Y=200 $D=22
M5 1 2 1 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=13220 $Y=200 $D=22
M6 1 2 1 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=15740 $Y=200 $D=22
M7 1 2 1 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=18260 $Y=200 $D=22
M8 1 2 1 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=20780 $Y=200 $D=22
M9 1 2 1 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=23300 $Y=200 $D=22
M10 1 2 1 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=25820 $Y=200 $D=22
M11 1 2 1 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=28340 $Y=200 $D=22
M12 1 2 1 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=30860 $Y=200 $D=22
M13 1 2 1 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=33380 $Y=200 $D=22
M14 1 2 1 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=35900 $Y=200 $D=22
M15 1 2 1 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=38420 $Y=200 $D=22
M16 1 2 1 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=40940 $Y=200 $D=22
M17 1 2 1 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=43460 $Y=200 $D=22
M18 1 2 1 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=45980 $Y=200 $D=22
M19 1 2 1 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=48500 $Y=200 $D=22
M20 1 2 1 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=51020 $Y=200 $D=22
M21 1 2 1 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=53540 $Y=200 $D=22
M22 1 2 1 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=56060 $Y=200 $D=22
M23 1 2 1 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=58580 $Y=200 $D=22
M24 1 2 1 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=61100 $Y=200 $D=22
M25 1 2 1 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=63620 $Y=200 $D=22
M26 1 2 1 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=66140 $Y=200 $D=22
M27 1 2 1 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=68660 $Y=200 $D=22
M28 1 2 1 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=71180 $Y=200 $D=22
M29 1 2 1 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=73700 $Y=200 $D=22
M30 1 2 1 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=76220 $Y=200 $D=22
M31 1 2 1 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=78740 $Y=200 $D=22
M32 1 2 1 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=81260 $Y=200 $D=22
M33 1 2 1 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=83780 $Y=200 $D=22
M34 1 2 1 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=86300 $Y=200 $D=22
M35 1 2 1 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=88820 $Y=200 $D=22
M36 1 2 1 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=91340 $Y=200 $D=22
M37 1 2 1 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=93860 $Y=200 $D=22
M38 1 2 1 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=96380 $Y=200 $D=22
M39 1 2 1 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=98900 $Y=200 $D=22
M40 1 2 1 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=101420 $Y=200 $D=22
M41 1 2 1 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=103940 $Y=200 $D=22
M42 1 2 1 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=106460 $Y=200 $D=22
M43 1 2 1 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=108980 $Y=200 $D=22
M44 1 2 1 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=111500 $Y=200 $D=22
M45 1 2 1 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=114020 $Y=200 $D=22
M46 1 2 1 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=116540 $Y=200 $D=22
M47 1 2 1 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=119060 $Y=200 $D=22
M48 1 2 1 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=121580 $Y=200 $D=22
M49 1 2 1 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=124100 $Y=200 $D=22
M50 1 2 1 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=126620 $Y=200 $D=22
M51 1 2 1 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=129140 $Y=200 $D=22
M52 1 2 1 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=131660 $Y=200 $D=22
M53 1 2 1 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=134180 $Y=200 $D=22
M54 1 2 1 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=136700 $Y=200 $D=22
M55 1 2 1 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=139220 $Y=200 $D=22
M56 1 2 1 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=141740 $Y=200 $D=22
M57 1 2 1 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=144260 $Y=200 $D=22
M58 1 2 1 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=146780 $Y=200 $D=22
M59 1 2 1 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=149300 $Y=200 $D=22
M60 1 2 1 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=151820 $Y=200 $D=22
M61 1 2 1 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=1.67141e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=154340 $Y=200 $D=22
.ENDS
***************************************
.SUBCKT cpoly_p_CDNS_5887047866536 1 2
** N=2 EP=2 IP=0 FDC=164
M0 1 2 1 cpoly_p w=6e-06 l=2e-06 c=8.0712e-14 as=1.68e-13 ad=7.488e-13 ps=1.44e-06 pd=1.13684e-06 sim_w=2.88e-06 m_per_maxw=2.08333 numb_sub_cont=4 nfing=1 $X=620 $Y=200 $D=21
M1 1 2 1 cpoly_p w=6e-06 l=2e-06 c=8.0712e-14 as=2.1408e-13 ad=7.488e-13 ps=1.44e-06 pd=1.13684e-06 sim_w=2.88e-06 m_per_maxw=2.08333 numb_sub_cont=4 nfing=1 $X=3140 $Y=200 $D=21
M2 1 2 1 cpoly_p w=6e-06 l=2e-06 c=8.0712e-14 as=2.1408e-13 ad=7.488e-13 ps=1.44e-06 pd=1.13684e-06 sim_w=2.88e-06 m_per_maxw=2.08333 numb_sub_cont=4 nfing=1 $X=5660 $Y=200 $D=21
M3 1 2 1 cpoly_p w=6e-06 l=2e-06 c=8.0712e-14 as=2.1408e-13 ad=7.488e-13 ps=1.44e-06 pd=1.13684e-06 sim_w=2.88e-06 m_per_maxw=2.08333 numb_sub_cont=4 nfing=1 $X=8180 $Y=200 $D=21
M4 1 2 1 cpoly_p w=6e-06 l=2e-06 c=8.0712e-14 as=2.1408e-13 ad=7.488e-13 ps=1.44e-06 pd=1.13684e-06 sim_w=2.88e-06 m_per_maxw=2.08333 numb_sub_cont=4 nfing=1 $X=10700 $Y=200 $D=21
M5 1 2 1 cpoly_p w=6e-06 l=2e-06 c=8.0712e-14 as=2.1408e-13 ad=7.488e-13 ps=1.44e-06 pd=1.13684e-06 sim_w=2.88e-06 m_per_maxw=2.08333 numb_sub_cont=4 nfing=1 $X=13220 $Y=200 $D=21
M6 1 2 1 cpoly_p w=6e-06 l=2e-06 c=8.0712e-14 as=2.1408e-13 ad=7.488e-13 ps=1.44e-06 pd=1.13684e-06 sim_w=2.88e-06 m_per_maxw=2.08333 numb_sub_cont=4 nfing=1 $X=15740 $Y=200 $D=21
M7 1 2 1 cpoly_p w=6e-06 l=2e-06 c=8.0712e-14 as=2.1408e-13 ad=7.488e-13 ps=1.44e-06 pd=1.13684e-06 sim_w=2.88e-06 m_per_maxw=2.08333 numb_sub_cont=4 nfing=1 $X=18260 $Y=200 $D=21
M8 1 2 1 cpoly_p w=6e-06 l=2e-06 c=8.0712e-14 as=2.1408e-13 ad=7.488e-13 ps=1.44e-06 pd=1.13684e-06 sim_w=2.88e-06 m_per_maxw=2.08333 numb_sub_cont=4 nfing=1 $X=20780 $Y=200 $D=21
M9 1 2 1 cpoly_p w=6e-06 l=2e-06 c=8.0712e-14 as=2.1408e-13 ad=7.488e-13 ps=1.44e-06 pd=1.13684e-06 sim_w=2.88e-06 m_per_maxw=2.08333 numb_sub_cont=4 nfing=1 $X=23300 $Y=200 $D=21
M10 1 2 1 cpoly_p w=6e-06 l=2e-06 c=8.0712e-14 as=2.1408e-13 ad=7.488e-13 ps=1.44e-06 pd=1.13684e-06 sim_w=2.88e-06 m_per_maxw=2.08333 numb_sub_cont=4 nfing=1 $X=25820 $Y=200 $D=21
M11 1 2 1 cpoly_p w=6e-06 l=2e-06 c=8.0712e-14 as=2.1408e-13 ad=7.488e-13 ps=1.44e-06 pd=1.13684e-06 sim_w=2.88e-06 m_per_maxw=2.08333 numb_sub_cont=4 nfing=1 $X=28340 $Y=200 $D=21
M12 1 2 1 cpoly_p w=6e-06 l=2e-06 c=8.0712e-14 as=2.1408e-13 ad=7.488e-13 ps=1.44e-06 pd=1.13684e-06 sim_w=2.88e-06 m_per_maxw=2.08333 numb_sub_cont=4 nfing=1 $X=30860 $Y=200 $D=21
M13 1 2 1 cpoly_p w=6e-06 l=2e-06 c=8.0712e-14 as=2.1408e-13 ad=7.488e-13 ps=1.44e-06 pd=1.13684e-06 sim_w=2.88e-06 m_per_maxw=2.08333 numb_sub_cont=4 nfing=1 $X=33380 $Y=200 $D=21
M14 1 2 1 cpoly_p w=6e-06 l=2e-06 c=8.0712e-14 as=2.1408e-13 ad=7.488e-13 ps=1.44e-06 pd=1.13684e-06 sim_w=2.88e-06 m_per_maxw=2.08333 numb_sub_cont=4 nfing=1 $X=35900 $Y=200 $D=21
M15 1 2 1 cpoly_p w=6e-06 l=2e-06 c=8.0712e-14 as=2.1408e-13 ad=7.488e-13 ps=1.44e-06 pd=1.13684e-06 sim_w=2.88e-06 m_per_maxw=2.08333 numb_sub_cont=4 nfing=1 $X=38420 $Y=200 $D=21
M16 1 2 1 cpoly_p w=6e-06 l=2e-06 c=8.0712e-14 as=2.1408e-13 ad=7.488e-13 ps=1.44e-06 pd=1.13684e-06 sim_w=2.88e-06 m_per_maxw=2.08333 numb_sub_cont=4 nfing=1 $X=40940 $Y=200 $D=21
M17 1 2 1 cpoly_p w=6e-06 l=2e-06 c=8.0712e-14 as=2.1408e-13 ad=7.488e-13 ps=1.44e-06 pd=1.13684e-06 sim_w=2.88e-06 m_per_maxw=2.08333 numb_sub_cont=4 nfing=1 $X=43460 $Y=200 $D=21
M18 1 2 1 cpoly_p w=6e-06 l=2e-06 c=8.0712e-14 as=2.1408e-13 ad=7.488e-13 ps=1.44e-06 pd=1.13684e-06 sim_w=2.88e-06 m_per_maxw=2.08333 numb_sub_cont=4 nfing=1 $X=45980 $Y=200 $D=21
M19 1 2 1 cpoly_p w=6e-06 l=2e-06 c=8.0712e-14 as=2.1408e-13 ad=7.488e-13 ps=1.44e-06 pd=1.13684e-06 sim_w=2.88e-06 m_per_maxw=2.08333 numb_sub_cont=4 nfing=1 $X=48500 $Y=200 $D=21
M20 1 2 1 cpoly_p w=6e-06 l=2e-06 c=8.0712e-14 as=2.1408e-13 ad=7.488e-13 ps=1.44e-06 pd=1.13684e-06 sim_w=2.88e-06 m_per_maxw=2.08333 numb_sub_cont=4 nfing=1 $X=51020 $Y=200 $D=21
M21 1 2 1 cpoly_p w=6e-06 l=2e-06 c=8.0712e-14 as=2.1408e-13 ad=7.488e-13 ps=1.44e-06 pd=1.13684e-06 sim_w=2.88e-06 m_per_maxw=2.08333 numb_sub_cont=4 nfing=1 $X=53540 $Y=200 $D=21
M22 1 2 1 cpoly_p w=6e-06 l=2e-06 c=8.0712e-14 as=2.1408e-13 ad=7.488e-13 ps=1.44e-06 pd=1.13684e-06 sim_w=2.88e-06 m_per_maxw=2.08333 numb_sub_cont=4 nfing=1 $X=56060 $Y=200 $D=21
M23 1 2 1 cpoly_p w=6e-06 l=2e-06 c=8.0712e-14 as=2.1408e-13 ad=7.488e-13 ps=1.44e-06 pd=1.13684e-06 sim_w=2.88e-06 m_per_maxw=2.08333 numb_sub_cont=4 nfing=1 $X=58580 $Y=200 $D=21
M24 1 2 1 cpoly_p w=6e-06 l=2e-06 c=8.0712e-14 as=2.1408e-13 ad=7.488e-13 ps=1.44e-06 pd=1.13684e-06 sim_w=2.88e-06 m_per_maxw=2.08333 numb_sub_cont=4 nfing=1 $X=61100 $Y=200 $D=21
M25 1 2 1 cpoly_p w=6e-06 l=2e-06 c=8.0712e-14 as=2.1408e-13 ad=7.488e-13 ps=1.44e-06 pd=1.13684e-06 sim_w=2.88e-06 m_per_maxw=2.08333 numb_sub_cont=4 nfing=1 $X=63620 $Y=200 $D=21
M26 1 2 1 cpoly_p w=6e-06 l=2e-06 c=8.0712e-14 as=2.1408e-13 ad=7.488e-13 ps=1.44e-06 pd=1.13684e-06 sim_w=2.88e-06 m_per_maxw=2.08333 numb_sub_cont=4 nfing=1 $X=66140 $Y=200 $D=21
M27 1 2 1 cpoly_p w=6e-06 l=2e-06 c=8.0712e-14 as=2.1408e-13 ad=7.488e-13 ps=1.44e-06 pd=1.13684e-06 sim_w=2.88e-06 m_per_maxw=2.08333 numb_sub_cont=4 nfing=1 $X=68660 $Y=200 $D=21
M28 1 2 1 cpoly_p w=6e-06 l=2e-06 c=8.0712e-14 as=2.1408e-13 ad=7.488e-13 ps=1.44e-06 pd=1.13684e-06 sim_w=2.88e-06 m_per_maxw=2.08333 numb_sub_cont=4 nfing=1 $X=71180 $Y=200 $D=21
M29 1 2 1 cpoly_p w=6e-06 l=2e-06 c=8.0712e-14 as=2.1408e-13 ad=7.488e-13 ps=1.44e-06 pd=1.13684e-06 sim_w=2.88e-06 m_per_maxw=2.08333 numb_sub_cont=4 nfing=1 $X=73700 $Y=200 $D=21
M30 1 2 1 cpoly_p w=6e-06 l=2e-06 c=8.0712e-14 as=2.1408e-13 ad=7.488e-13 ps=1.44e-06 pd=1.13684e-06 sim_w=2.88e-06 m_per_maxw=2.08333 numb_sub_cont=4 nfing=1 $X=76220 $Y=200 $D=21
M31 1 2 1 cpoly_p w=6e-06 l=2e-06 c=8.0712e-14 as=2.1408e-13 ad=7.488e-13 ps=1.44e-06 pd=1.13684e-06 sim_w=2.88e-06 m_per_maxw=2.08333 numb_sub_cont=4 nfing=1 $X=78740 $Y=200 $D=21
M32 1 2 1 cpoly_p w=6e-06 l=2e-06 c=8.0712e-14 as=2.1408e-13 ad=7.488e-13 ps=1.44e-06 pd=1.13684e-06 sim_w=2.88e-06 m_per_maxw=2.08333 numb_sub_cont=4 nfing=1 $X=81260 $Y=200 $D=21
M33 1 2 1 cpoly_p w=6e-06 l=2e-06 c=8.0712e-14 as=2.1408e-13 ad=7.488e-13 ps=1.44e-06 pd=1.13684e-06 sim_w=2.88e-06 m_per_maxw=2.08333 numb_sub_cont=4 nfing=1 $X=83780 $Y=200 $D=21
M34 1 2 1 cpoly_p w=6e-06 l=2e-06 c=8.0712e-14 as=2.1408e-13 ad=7.488e-13 ps=1.44e-06 pd=1.13684e-06 sim_w=2.88e-06 m_per_maxw=2.08333 numb_sub_cont=4 nfing=1 $X=86300 $Y=200 $D=21
M35 1 2 1 cpoly_p w=6e-06 l=2e-06 c=8.0712e-14 as=2.1408e-13 ad=7.488e-13 ps=1.44e-06 pd=1.13684e-06 sim_w=2.88e-06 m_per_maxw=2.08333 numb_sub_cont=4 nfing=1 $X=88820 $Y=200 $D=21
M36 1 2 1 cpoly_p w=6e-06 l=2e-06 c=8.0712e-14 as=2.1408e-13 ad=7.488e-13 ps=1.44e-06 pd=1.13684e-06 sim_w=2.88e-06 m_per_maxw=2.08333 numb_sub_cont=4 nfing=1 $X=91340 $Y=200 $D=21
M37 1 2 1 cpoly_p w=6e-06 l=2e-06 c=8.0712e-14 as=2.1408e-13 ad=7.488e-13 ps=1.44e-06 pd=1.13684e-06 sim_w=2.88e-06 m_per_maxw=2.08333 numb_sub_cont=4 nfing=1 $X=93860 $Y=200 $D=21
M38 1 2 1 cpoly_p w=6e-06 l=2e-06 c=8.0712e-14 as=2.1408e-13 ad=7.488e-13 ps=1.44e-06 pd=1.13684e-06 sim_w=2.88e-06 m_per_maxw=2.08333 numb_sub_cont=4 nfing=1 $X=96380 $Y=200 $D=21
M39 1 2 1 cpoly_p w=6e-06 l=2e-06 c=8.0712e-14 as=2.1408e-13 ad=7.488e-13 ps=1.44e-06 pd=1.13684e-06 sim_w=2.88e-06 m_per_maxw=2.08333 numb_sub_cont=4 nfing=1 $X=98900 $Y=200 $D=21
M40 1 2 1 cpoly_p w=6e-06 l=2e-06 c=8.0712e-14 as=2.1408e-13 ad=7.488e-13 ps=1.44e-06 pd=1.13684e-06 sim_w=2.88e-06 m_per_maxw=2.08333 numb_sub_cont=4 nfing=1 $X=101420 $Y=200 $D=21
M41 1 2 1 cpoly_p w=6e-06 l=2e-06 c=8.0712e-14 as=2.1408e-13 ad=7.488e-13 ps=1.44e-06 pd=1.13684e-06 sim_w=2.88e-06 m_per_maxw=2.08333 numb_sub_cont=4 nfing=1 $X=103940 $Y=200 $D=21
M42 1 2 1 cpoly_p w=6e-06 l=2e-06 c=8.0712e-14 as=2.1408e-13 ad=7.488e-13 ps=1.44e-06 pd=1.13684e-06 sim_w=2.88e-06 m_per_maxw=2.08333 numb_sub_cont=4 nfing=1 $X=106460 $Y=200 $D=21
M43 1 2 1 cpoly_p w=6e-06 l=2e-06 c=8.0712e-14 as=2.1408e-13 ad=7.488e-13 ps=1.44e-06 pd=1.13684e-06 sim_w=2.88e-06 m_per_maxw=2.08333 numb_sub_cont=4 nfing=1 $X=108980 $Y=200 $D=21
M44 1 2 1 cpoly_p w=6e-06 l=2e-06 c=8.0712e-14 as=2.1408e-13 ad=7.488e-13 ps=1.44e-06 pd=1.13684e-06 sim_w=2.88e-06 m_per_maxw=2.08333 numb_sub_cont=4 nfing=1 $X=111500 $Y=200 $D=21
M45 1 2 1 cpoly_p w=6e-06 l=2e-06 c=8.0712e-14 as=2.1408e-13 ad=7.488e-13 ps=1.44e-06 pd=1.13684e-06 sim_w=2.88e-06 m_per_maxw=2.08333 numb_sub_cont=4 nfing=1 $X=114020 $Y=200 $D=21
M46 1 2 1 cpoly_p w=6e-06 l=2e-06 c=8.0712e-14 as=2.1408e-13 ad=7.488e-13 ps=1.44e-06 pd=1.13684e-06 sim_w=2.88e-06 m_per_maxw=2.08333 numb_sub_cont=4 nfing=1 $X=116540 $Y=200 $D=21
M47 1 2 1 cpoly_p w=6e-06 l=2e-06 c=8.0712e-14 as=2.1408e-13 ad=7.488e-13 ps=1.44e-06 pd=1.13684e-06 sim_w=2.88e-06 m_per_maxw=2.08333 numb_sub_cont=4 nfing=1 $X=119060 $Y=200 $D=21
M48 1 2 1 cpoly_p w=6e-06 l=2e-06 c=8.0712e-14 as=2.1408e-13 ad=7.488e-13 ps=1.44e-06 pd=1.13684e-06 sim_w=2.88e-06 m_per_maxw=2.08333 numb_sub_cont=4 nfing=1 $X=121580 $Y=200 $D=21
M49 1 2 1 cpoly_p w=6e-06 l=2e-06 c=8.0712e-14 as=2.1408e-13 ad=7.488e-13 ps=1.44e-06 pd=1.13684e-06 sim_w=2.88e-06 m_per_maxw=2.08333 numb_sub_cont=4 nfing=1 $X=124100 $Y=200 $D=21
M50 1 2 1 cpoly_p w=6e-06 l=2e-06 c=8.0712e-14 as=2.1408e-13 ad=7.488e-13 ps=1.44e-06 pd=1.13684e-06 sim_w=2.88e-06 m_per_maxw=2.08333 numb_sub_cont=4 nfing=1 $X=126620 $Y=200 $D=21
M51 1 2 1 cpoly_p w=6e-06 l=2e-06 c=8.0712e-14 as=2.1408e-13 ad=7.488e-13 ps=1.44e-06 pd=1.13684e-06 sim_w=2.88e-06 m_per_maxw=2.08333 numb_sub_cont=4 nfing=1 $X=129140 $Y=200 $D=21
M52 1 2 1 cpoly_p w=6e-06 l=2e-06 c=8.0712e-14 as=2.1408e-13 ad=7.488e-13 ps=1.44e-06 pd=1.13684e-06 sim_w=2.88e-06 m_per_maxw=2.08333 numb_sub_cont=4 nfing=1 $X=131660 $Y=200 $D=21
M53 1 2 1 cpoly_p w=6e-06 l=2e-06 c=8.0712e-14 as=2.1408e-13 ad=7.488e-13 ps=1.44e-06 pd=1.13684e-06 sim_w=2.88e-06 m_per_maxw=2.08333 numb_sub_cont=4 nfing=1 $X=134180 $Y=200 $D=21
M54 1 2 1 cpoly_p w=6e-06 l=2e-06 c=8.0712e-14 as=2.1408e-13 ad=7.488e-13 ps=1.44e-06 pd=1.13684e-06 sim_w=2.88e-06 m_per_maxw=2.08333 numb_sub_cont=4 nfing=1 $X=136700 $Y=200 $D=21
M55 1 2 1 cpoly_p w=6e-06 l=2e-06 c=8.0712e-14 as=2.1408e-13 ad=7.488e-13 ps=1.44e-06 pd=1.13684e-06 sim_w=2.88e-06 m_per_maxw=2.08333 numb_sub_cont=4 nfing=1 $X=139220 $Y=200 $D=21
M56 1 2 1 cpoly_p w=6e-06 l=2e-06 c=8.0712e-14 as=2.1408e-13 ad=7.488e-13 ps=1.44e-06 pd=1.13684e-06 sim_w=2.88e-06 m_per_maxw=2.08333 numb_sub_cont=4 nfing=1 $X=141740 $Y=200 $D=21
M57 1 2 1 cpoly_p w=6e-06 l=2e-06 c=8.0712e-14 as=2.1408e-13 ad=7.488e-13 ps=1.44e-06 pd=1.13684e-06 sim_w=2.88e-06 m_per_maxw=2.08333 numb_sub_cont=4 nfing=1 $X=144260 $Y=200 $D=21
M58 1 2 1 cpoly_p w=6e-06 l=2e-06 c=8.0712e-14 as=2.1408e-13 ad=7.488e-13 ps=1.44e-06 pd=1.13684e-06 sim_w=2.88e-06 m_per_maxw=2.08333 numb_sub_cont=4 nfing=1 $X=146780 $Y=200 $D=21
M59 1 2 1 cpoly_p w=6e-06 l=2e-06 c=8.0712e-14 as=2.1408e-13 ad=7.488e-13 ps=1.44e-06 pd=1.13684e-06 sim_w=2.88e-06 m_per_maxw=2.08333 numb_sub_cont=4 nfing=1 $X=149300 $Y=200 $D=21
M60 1 2 1 cpoly_p w=6e-06 l=2e-06 c=8.0712e-14 as=2.1408e-13 ad=7.488e-13 ps=1.44e-06 pd=1.13684e-06 sim_w=2.88e-06 m_per_maxw=2.08333 numb_sub_cont=4 nfing=1 $X=151820 $Y=200 $D=21
M61 1 2 1 cpoly_p w=6e-06 l=2e-06 c=8.0712e-14 as=2.1408e-13 ad=7.488e-13 ps=1.44e-06 pd=1.13684e-06 sim_w=2.88e-06 m_per_maxw=2.08333 numb_sub_cont=4 nfing=1 $X=154340 $Y=200 $D=21
M62 1 2 1 cpoly_p w=6e-06 l=2e-06 c=8.0712e-14 as=2.1408e-13 ad=7.488e-13 ps=1.44e-06 pd=1.13684e-06 sim_w=2.88e-06 m_per_maxw=2.08333 numb_sub_cont=4 nfing=1 $X=156860 $Y=200 $D=21
M63 1 2 1 cpoly_p w=6e-06 l=2e-06 c=8.0712e-14 as=2.1408e-13 ad=7.488e-13 ps=1.44e-06 pd=1.13684e-06 sim_w=2.88e-06 m_per_maxw=2.08333 numb_sub_cont=4 nfing=1 $X=159380 $Y=200 $D=21
M64 1 2 1 cpoly_p w=6e-06 l=2e-06 c=8.0712e-14 as=2.1408e-13 ad=7.488e-13 ps=1.44e-06 pd=1.13684e-06 sim_w=2.88e-06 m_per_maxw=2.08333 numb_sub_cont=4 nfing=1 $X=161900 $Y=200 $D=21
M65 1 2 1 cpoly_p w=6e-06 l=2e-06 c=8.0712e-14 as=2.1408e-13 ad=7.488e-13 ps=1.44e-06 pd=1.13684e-06 sim_w=2.88e-06 m_per_maxw=2.08333 numb_sub_cont=4 nfing=1 $X=164420 $Y=200 $D=21
M66 1 2 1 cpoly_p w=6e-06 l=2e-06 c=8.0712e-14 as=2.1408e-13 ad=7.488e-13 ps=1.44e-06 pd=1.13684e-06 sim_w=2.88e-06 m_per_maxw=2.08333 numb_sub_cont=4 nfing=1 $X=166940 $Y=200 $D=21
M67 1 2 1 cpoly_p w=6e-06 l=2e-06 c=8.0712e-14 as=2.1408e-13 ad=7.488e-13 ps=1.44e-06 pd=1.13684e-06 sim_w=2.88e-06 m_per_maxw=2.08333 numb_sub_cont=4 nfing=1 $X=169460 $Y=200 $D=21
M68 1 2 1 cpoly_p w=6e-06 l=2e-06 c=8.0712e-14 as=2.1408e-13 ad=7.488e-13 ps=1.44e-06 pd=1.13684e-06 sim_w=2.88e-06 m_per_maxw=2.08333 numb_sub_cont=4 nfing=1 $X=171980 $Y=200 $D=21
M69 1 2 1 cpoly_p w=6e-06 l=2e-06 c=8.0712e-14 as=2.1408e-13 ad=7.488e-13 ps=1.44e-06 pd=1.13684e-06 sim_w=2.88e-06 m_per_maxw=2.08333 numb_sub_cont=4 nfing=1 $X=174500 $Y=200 $D=21
M70 1 2 1 cpoly_p w=6e-06 l=2e-06 c=8.0712e-14 as=2.1408e-13 ad=7.488e-13 ps=1.44e-06 pd=1.13684e-06 sim_w=2.88e-06 m_per_maxw=2.08333 numb_sub_cont=4 nfing=1 $X=177020 $Y=200 $D=21
M71 1 2 1 cpoly_p w=6e-06 l=2e-06 c=8.0712e-14 as=2.1408e-13 ad=7.488e-13 ps=1.44e-06 pd=1.13684e-06 sim_w=2.88e-06 m_per_maxw=2.08333 numb_sub_cont=4 nfing=1 $X=179540 $Y=200 $D=21
M72 1 2 1 cpoly_p w=6e-06 l=2e-06 c=8.0712e-14 as=2.1408e-13 ad=7.488e-13 ps=1.44e-06 pd=1.13684e-06 sim_w=2.88e-06 m_per_maxw=2.08333 numb_sub_cont=4 nfing=1 $X=182060 $Y=200 $D=21
M73 1 2 1 cpoly_p w=6e-06 l=2e-06 c=8.0712e-14 as=2.1408e-13 ad=7.488e-13 ps=1.44e-06 pd=1.13684e-06 sim_w=2.88e-06 m_per_maxw=2.08333 numb_sub_cont=4 nfing=1 $X=184580 $Y=200 $D=21
M74 1 2 1 cpoly_p w=6e-06 l=2e-06 c=8.0712e-14 as=2.1408e-13 ad=7.488e-13 ps=1.44e-06 pd=1.13684e-06 sim_w=2.88e-06 m_per_maxw=2.08333 numb_sub_cont=4 nfing=1 $X=187100 $Y=200 $D=21
M75 1 2 1 cpoly_p w=6e-06 l=2e-06 c=8.0712e-14 as=2.1408e-13 ad=7.488e-13 ps=1.44e-06 pd=1.13684e-06 sim_w=2.88e-06 m_per_maxw=2.08333 numb_sub_cont=4 nfing=1 $X=189620 $Y=200 $D=21
M76 1 2 1 cpoly_p w=6e-06 l=2e-06 c=8.0712e-14 as=2.1408e-13 ad=7.488e-13 ps=1.44e-06 pd=1.13684e-06 sim_w=2.88e-06 m_per_maxw=2.08333 numb_sub_cont=4 nfing=1 $X=192140 $Y=200 $D=21
M77 1 2 1 cpoly_p w=6e-06 l=2e-06 c=8.0712e-14 as=2.1408e-13 ad=7.488e-13 ps=1.44e-06 pd=1.13684e-06 sim_w=2.88e-06 m_per_maxw=2.08333 numb_sub_cont=4 nfing=1 $X=194660 $Y=200 $D=21
M78 1 2 1 cpoly_p w=6e-06 l=2e-06 c=8.0712e-14 as=2.1408e-13 ad=7.488e-13 ps=1.44e-06 pd=1.13684e-06 sim_w=2.88e-06 m_per_maxw=2.08333 numb_sub_cont=4 nfing=1 $X=197180 $Y=200 $D=21
M79 1 2 1 cpoly_p w=6e-06 l=2e-06 c=8.0712e-14 as=2.1408e-13 ad=7.488e-13 ps=1.44e-06 pd=1.13684e-06 sim_w=2.88e-06 m_per_maxw=2.08333 numb_sub_cont=4 nfing=1 $X=199700 $Y=200 $D=21
M80 1 2 1 cpoly_p w=6e-06 l=2e-06 c=8.0712e-14 as=2.1408e-13 ad=7.488e-13 ps=1.44e-06 pd=1.13684e-06 sim_w=2.88e-06 m_per_maxw=2.08333 numb_sub_cont=4 nfing=1 $X=202220 $Y=200 $D=21
M81 1 2 1 cpoly_p w=6e-06 l=2e-06 c=8.0712e-14 as=2.1408e-13 ad=7.488e-13 ps=1.44e-06 pd=1.13684e-06 sim_w=2.88e-06 m_per_maxw=2.08333 numb_sub_cont=4 nfing=1 $X=204740 $Y=200 $D=21
M82 1 2 1 cpoly_p w=6e-06 l=2e-06 c=8.0712e-14 as=2.1408e-13 ad=7.488e-13 ps=1.44e-06 pd=1.13684e-06 sim_w=2.88e-06 m_per_maxw=2.08333 numb_sub_cont=4 nfing=1 $X=207260 $Y=200 $D=21
M83 1 2 1 cpoly_p w=6e-06 l=2e-06 c=8.0712e-14 as=2.1408e-13 ad=7.488e-13 ps=1.44e-06 pd=1.13684e-06 sim_w=2.88e-06 m_per_maxw=2.08333 numb_sub_cont=4 nfing=1 $X=209780 $Y=200 $D=21
M84 1 2 1 cpoly_p w=6e-06 l=2e-06 c=8.0712e-14 as=2.1408e-13 ad=7.488e-13 ps=1.44e-06 pd=1.13684e-06 sim_w=2.88e-06 m_per_maxw=2.08333 numb_sub_cont=4 nfing=1 $X=212300 $Y=200 $D=21
M85 1 2 1 cpoly_p w=6e-06 l=2e-06 c=8.0712e-14 as=2.1408e-13 ad=7.488e-13 ps=1.44e-06 pd=1.13684e-06 sim_w=2.88e-06 m_per_maxw=2.08333 numb_sub_cont=4 nfing=1 $X=214820 $Y=200 $D=21
M86 1 2 1 cpoly_p w=6e-06 l=2e-06 c=8.0712e-14 as=2.1408e-13 ad=7.488e-13 ps=1.44e-06 pd=1.13684e-06 sim_w=2.88e-06 m_per_maxw=2.08333 numb_sub_cont=4 nfing=1 $X=217340 $Y=200 $D=21
M87 1 2 1 cpoly_p w=6e-06 l=2e-06 c=8.0712e-14 as=2.1408e-13 ad=7.488e-13 ps=1.44e-06 pd=1.13684e-06 sim_w=2.88e-06 m_per_maxw=2.08333 numb_sub_cont=4 nfing=1 $X=219860 $Y=200 $D=21
M88 1 2 1 cpoly_p w=6e-06 l=2e-06 c=8.0712e-14 as=2.1408e-13 ad=7.488e-13 ps=1.44e-06 pd=1.13684e-06 sim_w=2.88e-06 m_per_maxw=2.08333 numb_sub_cont=4 nfing=1 $X=222380 $Y=200 $D=21
M89 1 2 1 cpoly_p w=6e-06 l=2e-06 c=8.0712e-14 as=2.1408e-13 ad=7.488e-13 ps=1.44e-06 pd=1.13684e-06 sim_w=2.88e-06 m_per_maxw=2.08333 numb_sub_cont=4 nfing=1 $X=224900 $Y=200 $D=21
M90 1 2 1 cpoly_p w=6e-06 l=2e-06 c=8.0712e-14 as=2.1408e-13 ad=7.488e-13 ps=1.44e-06 pd=1.13684e-06 sim_w=2.88e-06 m_per_maxw=2.08333 numb_sub_cont=4 nfing=1 $X=227420 $Y=200 $D=21
M91 1 2 1 cpoly_p w=6e-06 l=2e-06 c=8.0712e-14 as=2.1408e-13 ad=7.488e-13 ps=1.44e-06 pd=1.13684e-06 sim_w=2.88e-06 m_per_maxw=2.08333 numb_sub_cont=4 nfing=1 $X=229940 $Y=200 $D=21
M92 1 2 1 cpoly_p w=6e-06 l=2e-06 c=8.0712e-14 as=2.1408e-13 ad=7.488e-13 ps=1.44e-06 pd=1.13684e-06 sim_w=2.88e-06 m_per_maxw=2.08333 numb_sub_cont=4 nfing=1 $X=232460 $Y=200 $D=21
M93 1 2 1 cpoly_p w=6e-06 l=2e-06 c=8.0712e-14 as=2.1408e-13 ad=7.488e-13 ps=1.44e-06 pd=1.13684e-06 sim_w=2.88e-06 m_per_maxw=2.08333 numb_sub_cont=4 nfing=1 $X=234980 $Y=200 $D=21
M94 1 2 1 cpoly_p w=6e-06 l=2e-06 c=8.0712e-14 as=2.1408e-13 ad=7.488e-13 ps=1.44e-06 pd=1.13684e-06 sim_w=2.88e-06 m_per_maxw=2.08333 numb_sub_cont=4 nfing=1 $X=237500 $Y=200 $D=21
M95 1 2 1 cpoly_p w=6e-06 l=2e-06 c=8.0712e-14 as=2.1408e-13 ad=7.488e-13 ps=1.44e-06 pd=1.13684e-06 sim_w=2.88e-06 m_per_maxw=2.08333 numb_sub_cont=4 nfing=1 $X=240020 $Y=200 $D=21
M96 1 2 1 cpoly_p w=6e-06 l=2e-06 c=8.0712e-14 as=2.1408e-13 ad=7.488e-13 ps=1.44e-06 pd=1.13684e-06 sim_w=2.88e-06 m_per_maxw=2.08333 numb_sub_cont=4 nfing=1 $X=242540 $Y=200 $D=21
M97 1 2 1 cpoly_p w=6e-06 l=2e-06 c=8.0712e-14 as=2.1408e-13 ad=7.488e-13 ps=1.44e-06 pd=1.13684e-06 sim_w=2.88e-06 m_per_maxw=2.08333 numb_sub_cont=4 nfing=1 $X=245060 $Y=200 $D=21
M98 1 2 1 cpoly_p w=6e-06 l=2e-06 c=8.0712e-14 as=2.1408e-13 ad=7.488e-13 ps=1.44e-06 pd=1.13684e-06 sim_w=2.88e-06 m_per_maxw=2.08333 numb_sub_cont=4 nfing=1 $X=247580 $Y=200 $D=21
M99 1 2 1 cpoly_p w=6e-06 l=2e-06 c=8.0712e-14 as=2.1408e-13 ad=7.488e-13 ps=1.44e-06 pd=1.13684e-06 sim_w=2.88e-06 m_per_maxw=2.08333 numb_sub_cont=4 nfing=1 $X=250100 $Y=200 $D=21
M100 1 2 1 cpoly_p w=6e-06 l=2e-06 c=8.0712e-14 as=2.1408e-13 ad=7.488e-13 ps=1.44e-06 pd=1.13684e-06 sim_w=2.88e-06 m_per_maxw=2.08333 numb_sub_cont=4 nfing=1 $X=252620 $Y=200 $D=21
M101 1 2 1 cpoly_p w=6e-06 l=2e-06 c=8.0712e-14 as=2.1408e-13 ad=7.488e-13 ps=1.44e-06 pd=1.13684e-06 sim_w=2.88e-06 m_per_maxw=2.08333 numb_sub_cont=4 nfing=1 $X=255140 $Y=200 $D=21
M102 1 2 1 cpoly_p w=6e-06 l=2e-06 c=8.0712e-14 as=2.1408e-13 ad=7.488e-13 ps=1.44e-06 pd=1.13684e-06 sim_w=2.88e-06 m_per_maxw=2.08333 numb_sub_cont=4 nfing=1 $X=257660 $Y=200 $D=21
M103 1 2 1 cpoly_p w=6e-06 l=2e-06 c=8.0712e-14 as=2.1408e-13 ad=7.488e-13 ps=1.44e-06 pd=1.13684e-06 sim_w=2.88e-06 m_per_maxw=2.08333 numb_sub_cont=4 nfing=1 $X=260180 $Y=200 $D=21
M104 1 2 1 cpoly_p w=6e-06 l=2e-06 c=8.0712e-14 as=2.1408e-13 ad=7.488e-13 ps=1.44e-06 pd=1.13684e-06 sim_w=2.88e-06 m_per_maxw=2.08333 numb_sub_cont=4 nfing=1 $X=262700 $Y=200 $D=21
M105 1 2 1 cpoly_p w=6e-06 l=2e-06 c=8.0712e-14 as=2.1408e-13 ad=7.488e-13 ps=1.44e-06 pd=1.13684e-06 sim_w=2.88e-06 m_per_maxw=2.08333 numb_sub_cont=4 nfing=1 $X=265220 $Y=200 $D=21
M106 1 2 1 cpoly_p w=6e-06 l=2e-06 c=8.0712e-14 as=2.1408e-13 ad=7.488e-13 ps=1.44e-06 pd=1.13684e-06 sim_w=2.88e-06 m_per_maxw=2.08333 numb_sub_cont=4 nfing=1 $X=267740 $Y=200 $D=21
M107 1 2 1 cpoly_p w=6e-06 l=2e-06 c=8.0712e-14 as=2.1408e-13 ad=7.488e-13 ps=1.44e-06 pd=1.13684e-06 sim_w=2.88e-06 m_per_maxw=2.08333 numb_sub_cont=4 nfing=1 $X=270260 $Y=200 $D=21
M108 1 2 1 cpoly_p w=6e-06 l=2e-06 c=8.0712e-14 as=2.1408e-13 ad=7.488e-13 ps=1.44e-06 pd=1.13684e-06 sim_w=2.88e-06 m_per_maxw=2.08333 numb_sub_cont=4 nfing=1 $X=272780 $Y=200 $D=21
M109 1 2 1 cpoly_p w=6e-06 l=2e-06 c=8.0712e-14 as=2.1408e-13 ad=7.488e-13 ps=1.44e-06 pd=1.13684e-06 sim_w=2.88e-06 m_per_maxw=2.08333 numb_sub_cont=4 nfing=1 $X=275300 $Y=200 $D=21
M110 1 2 1 cpoly_p w=6e-06 l=2e-06 c=8.0712e-14 as=2.1408e-13 ad=7.488e-13 ps=1.44e-06 pd=1.13684e-06 sim_w=2.88e-06 m_per_maxw=2.08333 numb_sub_cont=4 nfing=1 $X=277820 $Y=200 $D=21
M111 1 2 1 cpoly_p w=6e-06 l=2e-06 c=8.0712e-14 as=2.1408e-13 ad=7.488e-13 ps=1.44e-06 pd=1.13684e-06 sim_w=2.88e-06 m_per_maxw=2.08333 numb_sub_cont=4 nfing=1 $X=280340 $Y=200 $D=21
M112 1 2 1 cpoly_p w=6e-06 l=2e-06 c=8.0712e-14 as=2.1408e-13 ad=7.488e-13 ps=1.44e-06 pd=1.13684e-06 sim_w=2.88e-06 m_per_maxw=2.08333 numb_sub_cont=4 nfing=1 $X=282860 $Y=200 $D=21
M113 1 2 1 cpoly_p w=6e-06 l=2e-06 c=8.0712e-14 as=2.1408e-13 ad=7.488e-13 ps=1.44e-06 pd=1.13684e-06 sim_w=2.88e-06 m_per_maxw=2.08333 numb_sub_cont=4 nfing=1 $X=285380 $Y=200 $D=21
M114 1 2 1 cpoly_p w=6e-06 l=2e-06 c=8.0712e-14 as=2.1408e-13 ad=7.488e-13 ps=1.44e-06 pd=1.13684e-06 sim_w=2.88e-06 m_per_maxw=2.08333 numb_sub_cont=4 nfing=1 $X=287900 $Y=200 $D=21
M115 1 2 1 cpoly_p w=6e-06 l=2e-06 c=8.0712e-14 as=2.1408e-13 ad=7.488e-13 ps=1.44e-06 pd=1.13684e-06 sim_w=2.88e-06 m_per_maxw=2.08333 numb_sub_cont=4 nfing=1 $X=290420 $Y=200 $D=21
M116 1 2 1 cpoly_p w=6e-06 l=2e-06 c=8.0712e-14 as=2.1408e-13 ad=7.488e-13 ps=1.44e-06 pd=1.13684e-06 sim_w=2.88e-06 m_per_maxw=2.08333 numb_sub_cont=4 nfing=1 $X=292940 $Y=200 $D=21
M117 1 2 1 cpoly_p w=6e-06 l=2e-06 c=8.0712e-14 as=2.1408e-13 ad=7.488e-13 ps=1.44e-06 pd=1.13684e-06 sim_w=2.88e-06 m_per_maxw=2.08333 numb_sub_cont=4 nfing=1 $X=295460 $Y=200 $D=21
M118 1 2 1 cpoly_p w=6e-06 l=2e-06 c=8.0712e-14 as=2.1408e-13 ad=7.488e-13 ps=1.44e-06 pd=1.13684e-06 sim_w=2.88e-06 m_per_maxw=2.08333 numb_sub_cont=4 nfing=1 $X=297980 $Y=200 $D=21
M119 1 2 1 cpoly_p w=6e-06 l=2e-06 c=8.0712e-14 as=2.1408e-13 ad=7.488e-13 ps=1.44e-06 pd=1.13684e-06 sim_w=2.88e-06 m_per_maxw=2.08333 numb_sub_cont=4 nfing=1 $X=300500 $Y=200 $D=21
M120 1 2 1 cpoly_p w=6e-06 l=2e-06 c=8.0712e-14 as=2.1408e-13 ad=7.488e-13 ps=1.44e-06 pd=1.13684e-06 sim_w=2.88e-06 m_per_maxw=2.08333 numb_sub_cont=4 nfing=1 $X=303020 $Y=200 $D=21
M121 1 2 1 cpoly_p w=6e-06 l=2e-06 c=8.0712e-14 as=2.1408e-13 ad=7.488e-13 ps=1.44e-06 pd=1.13684e-06 sim_w=2.88e-06 m_per_maxw=2.08333 numb_sub_cont=4 nfing=1 $X=305540 $Y=200 $D=21
M122 1 2 1 cpoly_p w=6e-06 l=2e-06 c=8.0712e-14 as=2.1408e-13 ad=7.488e-13 ps=1.44e-06 pd=1.13684e-06 sim_w=2.88e-06 m_per_maxw=2.08333 numb_sub_cont=4 nfing=1 $X=308060 $Y=200 $D=21
M123 1 2 1 cpoly_p w=6e-06 l=2e-06 c=8.0712e-14 as=2.1408e-13 ad=7.488e-13 ps=1.44e-06 pd=1.13684e-06 sim_w=2.88e-06 m_per_maxw=2.08333 numb_sub_cont=4 nfing=1 $X=310580 $Y=200 $D=21
M124 1 2 1 cpoly_p w=6e-06 l=2e-06 c=8.0712e-14 as=2.1408e-13 ad=7.488e-13 ps=1.44e-06 pd=1.13684e-06 sim_w=2.88e-06 m_per_maxw=2.08333 numb_sub_cont=4 nfing=1 $X=313100 $Y=200 $D=21
M125 1 2 1 cpoly_p w=6e-06 l=2e-06 c=8.0712e-14 as=2.1408e-13 ad=7.488e-13 ps=1.44e-06 pd=1.13684e-06 sim_w=2.88e-06 m_per_maxw=2.08333 numb_sub_cont=4 nfing=1 $X=315620 $Y=200 $D=21
M126 1 2 1 cpoly_p w=6e-06 l=2e-06 c=8.0712e-14 as=2.1408e-13 ad=7.488e-13 ps=1.44e-06 pd=1.13684e-06 sim_w=2.88e-06 m_per_maxw=2.08333 numb_sub_cont=4 nfing=1 $X=318140 $Y=200 $D=21
M127 1 2 1 cpoly_p w=6e-06 l=2e-06 c=8.0712e-14 as=2.1408e-13 ad=7.488e-13 ps=1.44e-06 pd=1.13684e-06 sim_w=2.88e-06 m_per_maxw=2.08333 numb_sub_cont=4 nfing=1 $X=320660 $Y=200 $D=21
M128 1 2 1 cpoly_p w=6e-06 l=2e-06 c=8.0712e-14 as=2.1408e-13 ad=7.488e-13 ps=1.44e-06 pd=1.13684e-06 sim_w=2.88e-06 m_per_maxw=2.08333 numb_sub_cont=4 nfing=1 $X=323180 $Y=200 $D=21
M129 1 2 1 cpoly_p w=6e-06 l=2e-06 c=8.0712e-14 as=2.1408e-13 ad=7.488e-13 ps=1.44e-06 pd=1.13684e-06 sim_w=2.88e-06 m_per_maxw=2.08333 numb_sub_cont=4 nfing=1 $X=325700 $Y=200 $D=21
M130 1 2 1 cpoly_p w=6e-06 l=2e-06 c=8.0712e-14 as=2.1408e-13 ad=7.488e-13 ps=1.44e-06 pd=1.13684e-06 sim_w=2.88e-06 m_per_maxw=2.08333 numb_sub_cont=4 nfing=1 $X=328220 $Y=200 $D=21
M131 1 2 1 cpoly_p w=6e-06 l=2e-06 c=8.0712e-14 as=2.1408e-13 ad=7.488e-13 ps=1.44e-06 pd=1.13684e-06 sim_w=2.88e-06 m_per_maxw=2.08333 numb_sub_cont=4 nfing=1 $X=330740 $Y=200 $D=21
M132 1 2 1 cpoly_p w=6e-06 l=2e-06 c=8.0712e-14 as=2.1408e-13 ad=7.488e-13 ps=1.44e-06 pd=1.13684e-06 sim_w=2.88e-06 m_per_maxw=2.08333 numb_sub_cont=4 nfing=1 $X=333260 $Y=200 $D=21
M133 1 2 1 cpoly_p w=6e-06 l=2e-06 c=8.0712e-14 as=2.1408e-13 ad=7.488e-13 ps=1.44e-06 pd=1.13684e-06 sim_w=2.88e-06 m_per_maxw=2.08333 numb_sub_cont=4 nfing=1 $X=335780 $Y=200 $D=21
M134 1 2 1 cpoly_p w=6e-06 l=2e-06 c=8.0712e-14 as=2.1408e-13 ad=7.488e-13 ps=1.44e-06 pd=1.13684e-06 sim_w=2.88e-06 m_per_maxw=2.08333 numb_sub_cont=4 nfing=1 $X=338300 $Y=200 $D=21
M135 1 2 1 cpoly_p w=6e-06 l=2e-06 c=8.0712e-14 as=2.1408e-13 ad=7.488e-13 ps=1.44e-06 pd=1.13684e-06 sim_w=2.88e-06 m_per_maxw=2.08333 numb_sub_cont=4 nfing=1 $X=340820 $Y=200 $D=21
M136 1 2 1 cpoly_p w=6e-06 l=2e-06 c=8.0712e-14 as=2.1408e-13 ad=7.488e-13 ps=1.44e-06 pd=1.13684e-06 sim_w=2.88e-06 m_per_maxw=2.08333 numb_sub_cont=4 nfing=1 $X=343340 $Y=200 $D=21
M137 1 2 1 cpoly_p w=6e-06 l=2e-06 c=8.0712e-14 as=2.1408e-13 ad=7.488e-13 ps=1.44e-06 pd=1.13684e-06 sim_w=2.88e-06 m_per_maxw=2.08333 numb_sub_cont=4 nfing=1 $X=345860 $Y=200 $D=21
M138 1 2 1 cpoly_p w=6e-06 l=2e-06 c=8.0712e-14 as=2.1408e-13 ad=7.488e-13 ps=1.44e-06 pd=1.13684e-06 sim_w=2.88e-06 m_per_maxw=2.08333 numb_sub_cont=4 nfing=1 $X=348380 $Y=200 $D=21
M139 1 2 1 cpoly_p w=6e-06 l=2e-06 c=8.0712e-14 as=2.1408e-13 ad=7.488e-13 ps=1.44e-06 pd=1.13684e-06 sim_w=2.88e-06 m_per_maxw=2.08333 numb_sub_cont=4 nfing=1 $X=350900 $Y=200 $D=21
M140 1 2 1 cpoly_p w=6e-06 l=2e-06 c=8.0712e-14 as=2.1408e-13 ad=7.488e-13 ps=1.44e-06 pd=1.13684e-06 sim_w=2.88e-06 m_per_maxw=2.08333 numb_sub_cont=4 nfing=1 $X=353420 $Y=200 $D=21
M141 1 2 1 cpoly_p w=6e-06 l=2e-06 c=8.0712e-14 as=2.1408e-13 ad=7.488e-13 ps=1.44e-06 pd=1.13684e-06 sim_w=2.88e-06 m_per_maxw=2.08333 numb_sub_cont=4 nfing=1 $X=355940 $Y=200 $D=21
M142 1 2 1 cpoly_p w=6e-06 l=2e-06 c=8.0712e-14 as=2.1408e-13 ad=7.488e-13 ps=1.44e-06 pd=1.13684e-06 sim_w=2.88e-06 m_per_maxw=2.08333 numb_sub_cont=4 nfing=1 $X=358460 $Y=200 $D=21
M143 1 2 1 cpoly_p w=6e-06 l=2e-06 c=8.0712e-14 as=2.1408e-13 ad=7.488e-13 ps=1.44e-06 pd=1.13684e-06 sim_w=2.88e-06 m_per_maxw=2.08333 numb_sub_cont=4 nfing=1 $X=360980 $Y=200 $D=21
M144 1 2 1 cpoly_p w=6e-06 l=2e-06 c=8.0712e-14 as=2.1408e-13 ad=7.488e-13 ps=1.44e-06 pd=1.13684e-06 sim_w=2.88e-06 m_per_maxw=2.08333 numb_sub_cont=4 nfing=1 $X=363500 $Y=200 $D=21
M145 1 2 1 cpoly_p w=6e-06 l=2e-06 c=8.0712e-14 as=2.1408e-13 ad=7.488e-13 ps=1.44e-06 pd=1.13684e-06 sim_w=2.88e-06 m_per_maxw=2.08333 numb_sub_cont=4 nfing=1 $X=366020 $Y=200 $D=21
M146 1 2 1 cpoly_p w=6e-06 l=2e-06 c=8.0712e-14 as=2.1408e-13 ad=7.488e-13 ps=1.44e-06 pd=1.13684e-06 sim_w=2.88e-06 m_per_maxw=2.08333 numb_sub_cont=4 nfing=1 $X=368540 $Y=200 $D=21
M147 1 2 1 cpoly_p w=6e-06 l=2e-06 c=8.0712e-14 as=2.1408e-13 ad=7.488e-13 ps=1.44e-06 pd=1.13684e-06 sim_w=2.88e-06 m_per_maxw=2.08333 numb_sub_cont=4 nfing=1 $X=371060 $Y=200 $D=21
M148 1 2 1 cpoly_p w=6e-06 l=2e-06 c=8.0712e-14 as=2.1408e-13 ad=7.488e-13 ps=1.44e-06 pd=1.13684e-06 sim_w=2.88e-06 m_per_maxw=2.08333 numb_sub_cont=4 nfing=1 $X=373580 $Y=200 $D=21
M149 1 2 1 cpoly_p w=6e-06 l=2e-06 c=8.0712e-14 as=2.1408e-13 ad=7.488e-13 ps=1.44e-06 pd=1.13684e-06 sim_w=2.88e-06 m_per_maxw=2.08333 numb_sub_cont=4 nfing=1 $X=376100 $Y=200 $D=21
M150 1 2 1 cpoly_p w=6e-06 l=2e-06 c=8.0712e-14 as=2.1408e-13 ad=7.488e-13 ps=1.44e-06 pd=1.13684e-06 sim_w=2.88e-06 m_per_maxw=2.08333 numb_sub_cont=4 nfing=1 $X=378620 $Y=200 $D=21
M151 1 2 1 cpoly_p w=6e-06 l=2e-06 c=8.0712e-14 as=2.1408e-13 ad=7.488e-13 ps=1.44e-06 pd=1.13684e-06 sim_w=2.88e-06 m_per_maxw=2.08333 numb_sub_cont=4 nfing=1 $X=381140 $Y=200 $D=21
M152 1 2 1 cpoly_p w=6e-06 l=2e-06 c=8.0712e-14 as=2.1408e-13 ad=7.488e-13 ps=1.44e-06 pd=1.13684e-06 sim_w=2.88e-06 m_per_maxw=2.08333 numb_sub_cont=4 nfing=1 $X=383660 $Y=200 $D=21
M153 1 2 1 cpoly_p w=6e-06 l=2e-06 c=8.0712e-14 as=2.1408e-13 ad=7.488e-13 ps=1.44e-06 pd=1.13684e-06 sim_w=2.88e-06 m_per_maxw=2.08333 numb_sub_cont=4 nfing=1 $X=386180 $Y=200 $D=21
M154 1 2 1 cpoly_p w=6e-06 l=2e-06 c=8.0712e-14 as=2.1408e-13 ad=7.488e-13 ps=1.44e-06 pd=1.13684e-06 sim_w=2.88e-06 m_per_maxw=2.08333 numb_sub_cont=4 nfing=1 $X=388700 $Y=200 $D=21
M155 1 2 1 cpoly_p w=6e-06 l=2e-06 c=8.0712e-14 as=2.1408e-13 ad=7.488e-13 ps=1.44e-06 pd=1.13684e-06 sim_w=2.88e-06 m_per_maxw=2.08333 numb_sub_cont=4 nfing=1 $X=391220 $Y=200 $D=21
M156 1 2 1 cpoly_p w=6e-06 l=2e-06 c=8.0712e-14 as=2.1408e-13 ad=7.488e-13 ps=1.44e-06 pd=1.13684e-06 sim_w=2.88e-06 m_per_maxw=2.08333 numb_sub_cont=4 nfing=1 $X=393740 $Y=200 $D=21
M157 1 2 1 cpoly_p w=6e-06 l=2e-06 c=8.0712e-14 as=2.1408e-13 ad=7.488e-13 ps=1.44e-06 pd=1.13684e-06 sim_w=2.88e-06 m_per_maxw=2.08333 numb_sub_cont=4 nfing=1 $X=396260 $Y=200 $D=21
M158 1 2 1 cpoly_p w=6e-06 l=2e-06 c=8.0712e-14 as=2.1408e-13 ad=7.488e-13 ps=1.44e-06 pd=1.13684e-06 sim_w=2.88e-06 m_per_maxw=2.08333 numb_sub_cont=4 nfing=1 $X=398780 $Y=200 $D=21
M159 1 2 1 cpoly_p w=6e-06 l=2e-06 c=8.0712e-14 as=2.1408e-13 ad=7.488e-13 ps=1.44e-06 pd=1.13684e-06 sim_w=2.88e-06 m_per_maxw=2.08333 numb_sub_cont=4 nfing=1 $X=401300 $Y=200 $D=21
M160 1 2 1 cpoly_p w=6e-06 l=2e-06 c=8.0712e-14 as=2.1408e-13 ad=7.488e-13 ps=1.44e-06 pd=1.13684e-06 sim_w=2.88e-06 m_per_maxw=2.08333 numb_sub_cont=4 nfing=1 $X=403820 $Y=200 $D=21
M161 1 2 1 cpoly_p w=6e-06 l=2e-06 c=8.0712e-14 as=2.1408e-13 ad=7.488e-13 ps=1.44e-06 pd=1.13684e-06 sim_w=2.88e-06 m_per_maxw=2.08333 numb_sub_cont=4 nfing=1 $X=406340 $Y=200 $D=21
M162 1 2 1 cpoly_p w=6e-06 l=2e-06 c=8.0712e-14 as=2.1408e-13 ad=7.488e-13 ps=1.44e-06 pd=1.13684e-06 sim_w=2.88e-06 m_per_maxw=2.08333 numb_sub_cont=4 nfing=1 $X=408860 $Y=200 $D=21
M163 1 2 1 cpoly_p w=6e-06 l=2e-06 c=8.0712e-14 as=1.68e-13 ad=7.488e-13 ps=1.44e-06 pd=1.13684e-06 sim_w=2.88e-06 m_per_maxw=2.08333 numb_sub_cont=4 nfing=1 $X=411380 $Y=200 $D=21
.ENDS
***************************************
.SUBCKT cpoly_n_CDNS_5887047866529 1 2
** N=2 EP=2 IP=0 FDC=164
M0 1 2 1 cpoly_n w=6e-06 l=2e-06 c=7.5402e-14 as=2.4e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.4338e-06 sim_w=5.76e-06 m_per_maxw=1.04167 numb_sub_cont=3 nfing=1 $X=620 $Y=200 $D=22
M1 1 2 1 cpoly_n w=6e-06 l=2e-06 c=7.5402e-14 as=3.0336e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.4338e-06 sim_w=5.76e-06 m_per_maxw=1.04167 numb_sub_cont=3 nfing=1 $X=3140 $Y=200 $D=22
M2 1 2 1 cpoly_n w=6e-06 l=2e-06 c=7.5402e-14 as=3.0336e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.4338e-06 sim_w=5.76e-06 m_per_maxw=1.04167 numb_sub_cont=3 nfing=1 $X=5660 $Y=200 $D=22
M3 1 2 1 cpoly_n w=6e-06 l=2e-06 c=7.5402e-14 as=3.0336e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.4338e-06 sim_w=5.76e-06 m_per_maxw=1.04167 numb_sub_cont=3 nfing=1 $X=8180 $Y=200 $D=22
M4 1 2 1 cpoly_n w=6e-06 l=2e-06 c=7.5402e-14 as=3.0336e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.4338e-06 sim_w=5.76e-06 m_per_maxw=1.04167 numb_sub_cont=3 nfing=1 $X=10700 $Y=200 $D=22
M5 1 2 1 cpoly_n w=6e-06 l=2e-06 c=7.5402e-14 as=3.0336e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.4338e-06 sim_w=5.76e-06 m_per_maxw=1.04167 numb_sub_cont=3 nfing=1 $X=13220 $Y=200 $D=22
M6 1 2 1 cpoly_n w=6e-06 l=2e-06 c=7.5402e-14 as=3.0336e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.4338e-06 sim_w=5.76e-06 m_per_maxw=1.04167 numb_sub_cont=3 nfing=1 $X=15740 $Y=200 $D=22
M7 1 2 1 cpoly_n w=6e-06 l=2e-06 c=7.5402e-14 as=3.0336e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.4338e-06 sim_w=5.76e-06 m_per_maxw=1.04167 numb_sub_cont=3 nfing=1 $X=18260 $Y=200 $D=22
M8 1 2 1 cpoly_n w=6e-06 l=2e-06 c=7.5402e-14 as=3.0336e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.4338e-06 sim_w=5.76e-06 m_per_maxw=1.04167 numb_sub_cont=3 nfing=1 $X=20780 $Y=200 $D=22
M9 1 2 1 cpoly_n w=6e-06 l=2e-06 c=7.5402e-14 as=3.0336e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.4338e-06 sim_w=5.76e-06 m_per_maxw=1.04167 numb_sub_cont=3 nfing=1 $X=23300 $Y=200 $D=22
M10 1 2 1 cpoly_n w=6e-06 l=2e-06 c=7.5402e-14 as=3.0336e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.4338e-06 sim_w=5.76e-06 m_per_maxw=1.04167 numb_sub_cont=3 nfing=1 $X=25820 $Y=200 $D=22
M11 1 2 1 cpoly_n w=6e-06 l=2e-06 c=7.5402e-14 as=3.0336e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.4338e-06 sim_w=5.76e-06 m_per_maxw=1.04167 numb_sub_cont=3 nfing=1 $X=28340 $Y=200 $D=22
M12 1 2 1 cpoly_n w=6e-06 l=2e-06 c=7.5402e-14 as=3.0336e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.4338e-06 sim_w=5.76e-06 m_per_maxw=1.04167 numb_sub_cont=3 nfing=1 $X=30860 $Y=200 $D=22
M13 1 2 1 cpoly_n w=6e-06 l=2e-06 c=7.5402e-14 as=3.0336e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.4338e-06 sim_w=5.76e-06 m_per_maxw=1.04167 numb_sub_cont=3 nfing=1 $X=33380 $Y=200 $D=22
M14 1 2 1 cpoly_n w=6e-06 l=2e-06 c=7.5402e-14 as=3.0336e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.4338e-06 sim_w=5.76e-06 m_per_maxw=1.04167 numb_sub_cont=3 nfing=1 $X=35900 $Y=200 $D=22
M15 1 2 1 cpoly_n w=6e-06 l=2e-06 c=7.5402e-14 as=3.0336e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.4338e-06 sim_w=5.76e-06 m_per_maxw=1.04167 numb_sub_cont=3 nfing=1 $X=38420 $Y=200 $D=22
M16 1 2 1 cpoly_n w=6e-06 l=2e-06 c=7.5402e-14 as=3.0336e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.4338e-06 sim_w=5.76e-06 m_per_maxw=1.04167 numb_sub_cont=3 nfing=1 $X=40940 $Y=200 $D=22
M17 1 2 1 cpoly_n w=6e-06 l=2e-06 c=7.5402e-14 as=3.0336e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.4338e-06 sim_w=5.76e-06 m_per_maxw=1.04167 numb_sub_cont=3 nfing=1 $X=43460 $Y=200 $D=22
M18 1 2 1 cpoly_n w=6e-06 l=2e-06 c=7.5402e-14 as=3.0336e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.4338e-06 sim_w=5.76e-06 m_per_maxw=1.04167 numb_sub_cont=3 nfing=1 $X=45980 $Y=200 $D=22
M19 1 2 1 cpoly_n w=6e-06 l=2e-06 c=7.5402e-14 as=3.0336e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.4338e-06 sim_w=5.76e-06 m_per_maxw=1.04167 numb_sub_cont=3 nfing=1 $X=48500 $Y=200 $D=22
M20 1 2 1 cpoly_n w=6e-06 l=2e-06 c=7.5402e-14 as=3.0336e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.4338e-06 sim_w=5.76e-06 m_per_maxw=1.04167 numb_sub_cont=3 nfing=1 $X=51020 $Y=200 $D=22
M21 1 2 1 cpoly_n w=6e-06 l=2e-06 c=7.5402e-14 as=3.0336e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.4338e-06 sim_w=5.76e-06 m_per_maxw=1.04167 numb_sub_cont=3 nfing=1 $X=53540 $Y=200 $D=22
M22 1 2 1 cpoly_n w=6e-06 l=2e-06 c=7.5402e-14 as=3.0336e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.4338e-06 sim_w=5.76e-06 m_per_maxw=1.04167 numb_sub_cont=3 nfing=1 $X=56060 $Y=200 $D=22
M23 1 2 1 cpoly_n w=6e-06 l=2e-06 c=7.5402e-14 as=3.0336e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.4338e-06 sim_w=5.76e-06 m_per_maxw=1.04167 numb_sub_cont=3 nfing=1 $X=58580 $Y=200 $D=22
M24 1 2 1 cpoly_n w=6e-06 l=2e-06 c=7.5402e-14 as=3.0336e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.4338e-06 sim_w=5.76e-06 m_per_maxw=1.04167 numb_sub_cont=3 nfing=1 $X=61100 $Y=200 $D=22
M25 1 2 1 cpoly_n w=6e-06 l=2e-06 c=7.5402e-14 as=3.0336e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.4338e-06 sim_w=5.76e-06 m_per_maxw=1.04167 numb_sub_cont=3 nfing=1 $X=63620 $Y=200 $D=22
M26 1 2 1 cpoly_n w=6e-06 l=2e-06 c=7.5402e-14 as=3.0336e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.4338e-06 sim_w=5.76e-06 m_per_maxw=1.04167 numb_sub_cont=3 nfing=1 $X=66140 $Y=200 $D=22
M27 1 2 1 cpoly_n w=6e-06 l=2e-06 c=7.5402e-14 as=3.0336e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.4338e-06 sim_w=5.76e-06 m_per_maxw=1.04167 numb_sub_cont=3 nfing=1 $X=68660 $Y=200 $D=22
M28 1 2 1 cpoly_n w=6e-06 l=2e-06 c=7.5402e-14 as=3.0336e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.4338e-06 sim_w=5.76e-06 m_per_maxw=1.04167 numb_sub_cont=3 nfing=1 $X=71180 $Y=200 $D=22
M29 1 2 1 cpoly_n w=6e-06 l=2e-06 c=7.5402e-14 as=3.0336e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.4338e-06 sim_w=5.76e-06 m_per_maxw=1.04167 numb_sub_cont=3 nfing=1 $X=73700 $Y=200 $D=22
M30 1 2 1 cpoly_n w=6e-06 l=2e-06 c=7.5402e-14 as=3.0336e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.4338e-06 sim_w=5.76e-06 m_per_maxw=1.04167 numb_sub_cont=3 nfing=1 $X=76220 $Y=200 $D=22
M31 1 2 1 cpoly_n w=6e-06 l=2e-06 c=7.5402e-14 as=3.0336e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.4338e-06 sim_w=5.76e-06 m_per_maxw=1.04167 numb_sub_cont=3 nfing=1 $X=78740 $Y=200 $D=22
M32 1 2 1 cpoly_n w=6e-06 l=2e-06 c=7.5402e-14 as=3.0336e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.4338e-06 sim_w=5.76e-06 m_per_maxw=1.04167 numb_sub_cont=3 nfing=1 $X=81260 $Y=200 $D=22
M33 1 2 1 cpoly_n w=6e-06 l=2e-06 c=7.5402e-14 as=3.0336e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.4338e-06 sim_w=5.76e-06 m_per_maxw=1.04167 numb_sub_cont=3 nfing=1 $X=83780 $Y=200 $D=22
M34 1 2 1 cpoly_n w=6e-06 l=2e-06 c=7.5402e-14 as=3.0336e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.4338e-06 sim_w=5.76e-06 m_per_maxw=1.04167 numb_sub_cont=3 nfing=1 $X=86300 $Y=200 $D=22
M35 1 2 1 cpoly_n w=6e-06 l=2e-06 c=7.5402e-14 as=3.0336e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.4338e-06 sim_w=5.76e-06 m_per_maxw=1.04167 numb_sub_cont=3 nfing=1 $X=88820 $Y=200 $D=22
M36 1 2 1 cpoly_n w=6e-06 l=2e-06 c=7.5402e-14 as=3.0336e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.4338e-06 sim_w=5.76e-06 m_per_maxw=1.04167 numb_sub_cont=3 nfing=1 $X=91340 $Y=200 $D=22
M37 1 2 1 cpoly_n w=6e-06 l=2e-06 c=7.5402e-14 as=3.0336e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.4338e-06 sim_w=5.76e-06 m_per_maxw=1.04167 numb_sub_cont=3 nfing=1 $X=93860 $Y=200 $D=22
M38 1 2 1 cpoly_n w=6e-06 l=2e-06 c=7.5402e-14 as=3.0336e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.4338e-06 sim_w=5.76e-06 m_per_maxw=1.04167 numb_sub_cont=3 nfing=1 $X=96380 $Y=200 $D=22
M39 1 2 1 cpoly_n w=6e-06 l=2e-06 c=7.5402e-14 as=3.0336e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.4338e-06 sim_w=5.76e-06 m_per_maxw=1.04167 numb_sub_cont=3 nfing=1 $X=98900 $Y=200 $D=22
M40 1 2 1 cpoly_n w=6e-06 l=2e-06 c=7.5402e-14 as=3.0336e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.4338e-06 sim_w=5.76e-06 m_per_maxw=1.04167 numb_sub_cont=3 nfing=1 $X=101420 $Y=200 $D=22
M41 1 2 1 cpoly_n w=6e-06 l=2e-06 c=7.5402e-14 as=3.0336e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.4338e-06 sim_w=5.76e-06 m_per_maxw=1.04167 numb_sub_cont=3 nfing=1 $X=103940 $Y=200 $D=22
M42 1 2 1 cpoly_n w=6e-06 l=2e-06 c=7.5402e-14 as=3.0336e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.4338e-06 sim_w=5.76e-06 m_per_maxw=1.04167 numb_sub_cont=3 nfing=1 $X=106460 $Y=200 $D=22
M43 1 2 1 cpoly_n w=6e-06 l=2e-06 c=7.5402e-14 as=3.0336e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.4338e-06 sim_w=5.76e-06 m_per_maxw=1.04167 numb_sub_cont=3 nfing=1 $X=108980 $Y=200 $D=22
M44 1 2 1 cpoly_n w=6e-06 l=2e-06 c=7.5402e-14 as=3.0336e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.4338e-06 sim_w=5.76e-06 m_per_maxw=1.04167 numb_sub_cont=3 nfing=1 $X=111500 $Y=200 $D=22
M45 1 2 1 cpoly_n w=6e-06 l=2e-06 c=7.5402e-14 as=3.0336e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.4338e-06 sim_w=5.76e-06 m_per_maxw=1.04167 numb_sub_cont=3 nfing=1 $X=114020 $Y=200 $D=22
M46 1 2 1 cpoly_n w=6e-06 l=2e-06 c=7.5402e-14 as=3.0336e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.4338e-06 sim_w=5.76e-06 m_per_maxw=1.04167 numb_sub_cont=3 nfing=1 $X=116540 $Y=200 $D=22
M47 1 2 1 cpoly_n w=6e-06 l=2e-06 c=7.5402e-14 as=3.0336e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.4338e-06 sim_w=5.76e-06 m_per_maxw=1.04167 numb_sub_cont=3 nfing=1 $X=119060 $Y=200 $D=22
M48 1 2 1 cpoly_n w=6e-06 l=2e-06 c=7.5402e-14 as=3.0336e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.4338e-06 sim_w=5.76e-06 m_per_maxw=1.04167 numb_sub_cont=3 nfing=1 $X=121580 $Y=200 $D=22
M49 1 2 1 cpoly_n w=6e-06 l=2e-06 c=7.5402e-14 as=3.0336e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.4338e-06 sim_w=5.76e-06 m_per_maxw=1.04167 numb_sub_cont=3 nfing=1 $X=124100 $Y=200 $D=22
M50 1 2 1 cpoly_n w=6e-06 l=2e-06 c=7.5402e-14 as=3.0336e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.4338e-06 sim_w=5.76e-06 m_per_maxw=1.04167 numb_sub_cont=3 nfing=1 $X=126620 $Y=200 $D=22
M51 1 2 1 cpoly_n w=6e-06 l=2e-06 c=7.5402e-14 as=3.0336e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.4338e-06 sim_w=5.76e-06 m_per_maxw=1.04167 numb_sub_cont=3 nfing=1 $X=129140 $Y=200 $D=22
M52 1 2 1 cpoly_n w=6e-06 l=2e-06 c=7.5402e-14 as=3.0336e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.4338e-06 sim_w=5.76e-06 m_per_maxw=1.04167 numb_sub_cont=3 nfing=1 $X=131660 $Y=200 $D=22
M53 1 2 1 cpoly_n w=6e-06 l=2e-06 c=7.5402e-14 as=3.0336e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.4338e-06 sim_w=5.76e-06 m_per_maxw=1.04167 numb_sub_cont=3 nfing=1 $X=134180 $Y=200 $D=22
M54 1 2 1 cpoly_n w=6e-06 l=2e-06 c=7.5402e-14 as=3.0336e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.4338e-06 sim_w=5.76e-06 m_per_maxw=1.04167 numb_sub_cont=3 nfing=1 $X=136700 $Y=200 $D=22
M55 1 2 1 cpoly_n w=6e-06 l=2e-06 c=7.5402e-14 as=3.0336e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.4338e-06 sim_w=5.76e-06 m_per_maxw=1.04167 numb_sub_cont=3 nfing=1 $X=139220 $Y=200 $D=22
M56 1 2 1 cpoly_n w=6e-06 l=2e-06 c=7.5402e-14 as=3.0336e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.4338e-06 sim_w=5.76e-06 m_per_maxw=1.04167 numb_sub_cont=3 nfing=1 $X=141740 $Y=200 $D=22
M57 1 2 1 cpoly_n w=6e-06 l=2e-06 c=7.5402e-14 as=3.0336e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.4338e-06 sim_w=5.76e-06 m_per_maxw=1.04167 numb_sub_cont=3 nfing=1 $X=144260 $Y=200 $D=22
M58 1 2 1 cpoly_n w=6e-06 l=2e-06 c=7.5402e-14 as=3.0336e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.4338e-06 sim_w=5.76e-06 m_per_maxw=1.04167 numb_sub_cont=3 nfing=1 $X=146780 $Y=200 $D=22
M59 1 2 1 cpoly_n w=6e-06 l=2e-06 c=7.5402e-14 as=3.0336e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.4338e-06 sim_w=5.76e-06 m_per_maxw=1.04167 numb_sub_cont=3 nfing=1 $X=149300 $Y=200 $D=22
M60 1 2 1 cpoly_n w=6e-06 l=2e-06 c=7.5402e-14 as=3.0336e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.4338e-06 sim_w=5.76e-06 m_per_maxw=1.04167 numb_sub_cont=3 nfing=1 $X=151820 $Y=200 $D=22
M61 1 2 1 cpoly_n w=6e-06 l=2e-06 c=7.5402e-14 as=3.0336e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.4338e-06 sim_w=5.76e-06 m_per_maxw=1.04167 numb_sub_cont=3 nfing=1 $X=154340 $Y=200 $D=22
M62 1 2 1 cpoly_n w=6e-06 l=2e-06 c=7.5402e-14 as=3.0336e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.4338e-06 sim_w=5.76e-06 m_per_maxw=1.04167 numb_sub_cont=3 nfing=1 $X=156860 $Y=200 $D=22
M63 1 2 1 cpoly_n w=6e-06 l=2e-06 c=7.5402e-14 as=3.0336e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.4338e-06 sim_w=5.76e-06 m_per_maxw=1.04167 numb_sub_cont=3 nfing=1 $X=159380 $Y=200 $D=22
M64 1 2 1 cpoly_n w=6e-06 l=2e-06 c=7.5402e-14 as=3.0336e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.4338e-06 sim_w=5.76e-06 m_per_maxw=1.04167 numb_sub_cont=3 nfing=1 $X=161900 $Y=200 $D=22
M65 1 2 1 cpoly_n w=6e-06 l=2e-06 c=7.5402e-14 as=3.0336e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.4338e-06 sim_w=5.76e-06 m_per_maxw=1.04167 numb_sub_cont=3 nfing=1 $X=164420 $Y=200 $D=22
M66 1 2 1 cpoly_n w=6e-06 l=2e-06 c=7.5402e-14 as=3.0336e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.4338e-06 sim_w=5.76e-06 m_per_maxw=1.04167 numb_sub_cont=3 nfing=1 $X=166940 $Y=200 $D=22
M67 1 2 1 cpoly_n w=6e-06 l=2e-06 c=7.5402e-14 as=3.0336e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.4338e-06 sim_w=5.76e-06 m_per_maxw=1.04167 numb_sub_cont=3 nfing=1 $X=169460 $Y=200 $D=22
M68 1 2 1 cpoly_n w=6e-06 l=2e-06 c=7.5402e-14 as=3.0336e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.4338e-06 sim_w=5.76e-06 m_per_maxw=1.04167 numb_sub_cont=3 nfing=1 $X=171980 $Y=200 $D=22
M69 1 2 1 cpoly_n w=6e-06 l=2e-06 c=7.5402e-14 as=3.0336e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.4338e-06 sim_w=5.76e-06 m_per_maxw=1.04167 numb_sub_cont=3 nfing=1 $X=174500 $Y=200 $D=22
M70 1 2 1 cpoly_n w=6e-06 l=2e-06 c=7.5402e-14 as=3.0336e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.4338e-06 sim_w=5.76e-06 m_per_maxw=1.04167 numb_sub_cont=3 nfing=1 $X=177020 $Y=200 $D=22
M71 1 2 1 cpoly_n w=6e-06 l=2e-06 c=7.5402e-14 as=3.0336e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.4338e-06 sim_w=5.76e-06 m_per_maxw=1.04167 numb_sub_cont=3 nfing=1 $X=179540 $Y=200 $D=22
M72 1 2 1 cpoly_n w=6e-06 l=2e-06 c=7.5402e-14 as=3.0336e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.4338e-06 sim_w=5.76e-06 m_per_maxw=1.04167 numb_sub_cont=3 nfing=1 $X=182060 $Y=200 $D=22
M73 1 2 1 cpoly_n w=6e-06 l=2e-06 c=7.5402e-14 as=3.0336e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.4338e-06 sim_w=5.76e-06 m_per_maxw=1.04167 numb_sub_cont=3 nfing=1 $X=184580 $Y=200 $D=22
M74 1 2 1 cpoly_n w=6e-06 l=2e-06 c=7.5402e-14 as=3.0336e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.4338e-06 sim_w=5.76e-06 m_per_maxw=1.04167 numb_sub_cont=3 nfing=1 $X=187100 $Y=200 $D=22
M75 1 2 1 cpoly_n w=6e-06 l=2e-06 c=7.5402e-14 as=3.0336e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.4338e-06 sim_w=5.76e-06 m_per_maxw=1.04167 numb_sub_cont=3 nfing=1 $X=189620 $Y=200 $D=22
M76 1 2 1 cpoly_n w=6e-06 l=2e-06 c=7.5402e-14 as=3.0336e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.4338e-06 sim_w=5.76e-06 m_per_maxw=1.04167 numb_sub_cont=3 nfing=1 $X=192140 $Y=200 $D=22
M77 1 2 1 cpoly_n w=6e-06 l=2e-06 c=7.5402e-14 as=3.0336e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.4338e-06 sim_w=5.76e-06 m_per_maxw=1.04167 numb_sub_cont=3 nfing=1 $X=194660 $Y=200 $D=22
M78 1 2 1 cpoly_n w=6e-06 l=2e-06 c=7.5402e-14 as=3.0336e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.4338e-06 sim_w=5.76e-06 m_per_maxw=1.04167 numb_sub_cont=3 nfing=1 $X=197180 $Y=200 $D=22
M79 1 2 1 cpoly_n w=6e-06 l=2e-06 c=7.5402e-14 as=3.0336e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.4338e-06 sim_w=5.76e-06 m_per_maxw=1.04167 numb_sub_cont=3 nfing=1 $X=199700 $Y=200 $D=22
M80 1 2 1 cpoly_n w=6e-06 l=2e-06 c=7.5402e-14 as=3.0336e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.4338e-06 sim_w=5.76e-06 m_per_maxw=1.04167 numb_sub_cont=3 nfing=1 $X=202220 $Y=200 $D=22
M81 1 2 1 cpoly_n w=6e-06 l=2e-06 c=7.5402e-14 as=3.0336e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.4338e-06 sim_w=5.76e-06 m_per_maxw=1.04167 numb_sub_cont=3 nfing=1 $X=204740 $Y=200 $D=22
M82 1 2 1 cpoly_n w=6e-06 l=2e-06 c=7.5402e-14 as=3.0336e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.4338e-06 sim_w=5.76e-06 m_per_maxw=1.04167 numb_sub_cont=3 nfing=1 $X=207260 $Y=200 $D=22
M83 1 2 1 cpoly_n w=6e-06 l=2e-06 c=7.5402e-14 as=3.0336e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.4338e-06 sim_w=5.76e-06 m_per_maxw=1.04167 numb_sub_cont=3 nfing=1 $X=209780 $Y=200 $D=22
M84 1 2 1 cpoly_n w=6e-06 l=2e-06 c=7.5402e-14 as=3.0336e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.4338e-06 sim_w=5.76e-06 m_per_maxw=1.04167 numb_sub_cont=3 nfing=1 $X=212300 $Y=200 $D=22
M85 1 2 1 cpoly_n w=6e-06 l=2e-06 c=7.5402e-14 as=3.0336e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.4338e-06 sim_w=5.76e-06 m_per_maxw=1.04167 numb_sub_cont=3 nfing=1 $X=214820 $Y=200 $D=22
M86 1 2 1 cpoly_n w=6e-06 l=2e-06 c=7.5402e-14 as=3.0336e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.4338e-06 sim_w=5.76e-06 m_per_maxw=1.04167 numb_sub_cont=3 nfing=1 $X=217340 $Y=200 $D=22
M87 1 2 1 cpoly_n w=6e-06 l=2e-06 c=7.5402e-14 as=3.0336e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.4338e-06 sim_w=5.76e-06 m_per_maxw=1.04167 numb_sub_cont=3 nfing=1 $X=219860 $Y=200 $D=22
M88 1 2 1 cpoly_n w=6e-06 l=2e-06 c=7.5402e-14 as=3.0336e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.4338e-06 sim_w=5.76e-06 m_per_maxw=1.04167 numb_sub_cont=3 nfing=1 $X=222380 $Y=200 $D=22
M89 1 2 1 cpoly_n w=6e-06 l=2e-06 c=7.5402e-14 as=3.0336e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.4338e-06 sim_w=5.76e-06 m_per_maxw=1.04167 numb_sub_cont=3 nfing=1 $X=224900 $Y=200 $D=22
M90 1 2 1 cpoly_n w=6e-06 l=2e-06 c=7.5402e-14 as=3.0336e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.4338e-06 sim_w=5.76e-06 m_per_maxw=1.04167 numb_sub_cont=3 nfing=1 $X=227420 $Y=200 $D=22
M91 1 2 1 cpoly_n w=6e-06 l=2e-06 c=7.5402e-14 as=3.0336e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.4338e-06 sim_w=5.76e-06 m_per_maxw=1.04167 numb_sub_cont=3 nfing=1 $X=229940 $Y=200 $D=22
M92 1 2 1 cpoly_n w=6e-06 l=2e-06 c=7.5402e-14 as=3.0336e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.4338e-06 sim_w=5.76e-06 m_per_maxw=1.04167 numb_sub_cont=3 nfing=1 $X=232460 $Y=200 $D=22
M93 1 2 1 cpoly_n w=6e-06 l=2e-06 c=7.5402e-14 as=3.0336e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.4338e-06 sim_w=5.76e-06 m_per_maxw=1.04167 numb_sub_cont=3 nfing=1 $X=234980 $Y=200 $D=22
M94 1 2 1 cpoly_n w=6e-06 l=2e-06 c=7.5402e-14 as=3.0336e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.4338e-06 sim_w=5.76e-06 m_per_maxw=1.04167 numb_sub_cont=3 nfing=1 $X=237500 $Y=200 $D=22
M95 1 2 1 cpoly_n w=6e-06 l=2e-06 c=7.5402e-14 as=3.0336e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.4338e-06 sim_w=5.76e-06 m_per_maxw=1.04167 numb_sub_cont=3 nfing=1 $X=240020 $Y=200 $D=22
M96 1 2 1 cpoly_n w=6e-06 l=2e-06 c=7.5402e-14 as=3.0336e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.4338e-06 sim_w=5.76e-06 m_per_maxw=1.04167 numb_sub_cont=3 nfing=1 $X=242540 $Y=200 $D=22
M97 1 2 1 cpoly_n w=6e-06 l=2e-06 c=7.5402e-14 as=3.0336e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.4338e-06 sim_w=5.76e-06 m_per_maxw=1.04167 numb_sub_cont=3 nfing=1 $X=245060 $Y=200 $D=22
M98 1 2 1 cpoly_n w=6e-06 l=2e-06 c=7.5402e-14 as=3.0336e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.4338e-06 sim_w=5.76e-06 m_per_maxw=1.04167 numb_sub_cont=3 nfing=1 $X=247580 $Y=200 $D=22
M99 1 2 1 cpoly_n w=6e-06 l=2e-06 c=7.5402e-14 as=3.0336e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.4338e-06 sim_w=5.76e-06 m_per_maxw=1.04167 numb_sub_cont=3 nfing=1 $X=250100 $Y=200 $D=22
M100 1 2 1 cpoly_n w=6e-06 l=2e-06 c=7.5402e-14 as=3.0336e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.4338e-06 sim_w=5.76e-06 m_per_maxw=1.04167 numb_sub_cont=3 nfing=1 $X=252620 $Y=200 $D=22
M101 1 2 1 cpoly_n w=6e-06 l=2e-06 c=7.5402e-14 as=3.0336e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.4338e-06 sim_w=5.76e-06 m_per_maxw=1.04167 numb_sub_cont=3 nfing=1 $X=255140 $Y=200 $D=22
M102 1 2 1 cpoly_n w=6e-06 l=2e-06 c=7.5402e-14 as=3.0336e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.4338e-06 sim_w=5.76e-06 m_per_maxw=1.04167 numb_sub_cont=3 nfing=1 $X=257660 $Y=200 $D=22
M103 1 2 1 cpoly_n w=6e-06 l=2e-06 c=7.5402e-14 as=3.0336e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.4338e-06 sim_w=5.76e-06 m_per_maxw=1.04167 numb_sub_cont=3 nfing=1 $X=260180 $Y=200 $D=22
M104 1 2 1 cpoly_n w=6e-06 l=2e-06 c=7.5402e-14 as=3.0336e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.4338e-06 sim_w=5.76e-06 m_per_maxw=1.04167 numb_sub_cont=3 nfing=1 $X=262700 $Y=200 $D=22
M105 1 2 1 cpoly_n w=6e-06 l=2e-06 c=7.5402e-14 as=3.0336e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.4338e-06 sim_w=5.76e-06 m_per_maxw=1.04167 numb_sub_cont=3 nfing=1 $X=265220 $Y=200 $D=22
M106 1 2 1 cpoly_n w=6e-06 l=2e-06 c=7.5402e-14 as=3.0336e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.4338e-06 sim_w=5.76e-06 m_per_maxw=1.04167 numb_sub_cont=3 nfing=1 $X=267740 $Y=200 $D=22
M107 1 2 1 cpoly_n w=6e-06 l=2e-06 c=7.5402e-14 as=3.0336e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.4338e-06 sim_w=5.76e-06 m_per_maxw=1.04167 numb_sub_cont=3 nfing=1 $X=270260 $Y=200 $D=22
M108 1 2 1 cpoly_n w=6e-06 l=2e-06 c=7.5402e-14 as=3.0336e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.4338e-06 sim_w=5.76e-06 m_per_maxw=1.04167 numb_sub_cont=3 nfing=1 $X=272780 $Y=200 $D=22
M109 1 2 1 cpoly_n w=6e-06 l=2e-06 c=7.5402e-14 as=3.0336e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.4338e-06 sim_w=5.76e-06 m_per_maxw=1.04167 numb_sub_cont=3 nfing=1 $X=275300 $Y=200 $D=22
M110 1 2 1 cpoly_n w=6e-06 l=2e-06 c=7.5402e-14 as=3.0336e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.4338e-06 sim_w=5.76e-06 m_per_maxw=1.04167 numb_sub_cont=3 nfing=1 $X=277820 $Y=200 $D=22
M111 1 2 1 cpoly_n w=6e-06 l=2e-06 c=7.5402e-14 as=3.0336e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.4338e-06 sim_w=5.76e-06 m_per_maxw=1.04167 numb_sub_cont=3 nfing=1 $X=280340 $Y=200 $D=22
M112 1 2 1 cpoly_n w=6e-06 l=2e-06 c=7.5402e-14 as=3.0336e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.4338e-06 sim_w=5.76e-06 m_per_maxw=1.04167 numb_sub_cont=3 nfing=1 $X=282860 $Y=200 $D=22
M113 1 2 1 cpoly_n w=6e-06 l=2e-06 c=7.5402e-14 as=3.0336e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.4338e-06 sim_w=5.76e-06 m_per_maxw=1.04167 numb_sub_cont=3 nfing=1 $X=285380 $Y=200 $D=22
M114 1 2 1 cpoly_n w=6e-06 l=2e-06 c=7.5402e-14 as=3.0336e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.4338e-06 sim_w=5.76e-06 m_per_maxw=1.04167 numb_sub_cont=3 nfing=1 $X=287900 $Y=200 $D=22
M115 1 2 1 cpoly_n w=6e-06 l=2e-06 c=7.5402e-14 as=3.0336e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.4338e-06 sim_w=5.76e-06 m_per_maxw=1.04167 numb_sub_cont=3 nfing=1 $X=290420 $Y=200 $D=22
M116 1 2 1 cpoly_n w=6e-06 l=2e-06 c=7.5402e-14 as=3.0336e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.4338e-06 sim_w=5.76e-06 m_per_maxw=1.04167 numb_sub_cont=3 nfing=1 $X=292940 $Y=200 $D=22
M117 1 2 1 cpoly_n w=6e-06 l=2e-06 c=7.5402e-14 as=3.0336e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.4338e-06 sim_w=5.76e-06 m_per_maxw=1.04167 numb_sub_cont=3 nfing=1 $X=295460 $Y=200 $D=22
M118 1 2 1 cpoly_n w=6e-06 l=2e-06 c=7.5402e-14 as=3.0336e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.4338e-06 sim_w=5.76e-06 m_per_maxw=1.04167 numb_sub_cont=3 nfing=1 $X=297980 $Y=200 $D=22
M119 1 2 1 cpoly_n w=6e-06 l=2e-06 c=7.5402e-14 as=3.0336e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.4338e-06 sim_w=5.76e-06 m_per_maxw=1.04167 numb_sub_cont=3 nfing=1 $X=300500 $Y=200 $D=22
M120 1 2 1 cpoly_n w=6e-06 l=2e-06 c=7.5402e-14 as=3.0336e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.4338e-06 sim_w=5.76e-06 m_per_maxw=1.04167 numb_sub_cont=3 nfing=1 $X=303020 $Y=200 $D=22
M121 1 2 1 cpoly_n w=6e-06 l=2e-06 c=7.5402e-14 as=3.0336e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.4338e-06 sim_w=5.76e-06 m_per_maxw=1.04167 numb_sub_cont=3 nfing=1 $X=305540 $Y=200 $D=22
M122 1 2 1 cpoly_n w=6e-06 l=2e-06 c=7.5402e-14 as=3.0336e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.4338e-06 sim_w=5.76e-06 m_per_maxw=1.04167 numb_sub_cont=3 nfing=1 $X=308060 $Y=200 $D=22
M123 1 2 1 cpoly_n w=6e-06 l=2e-06 c=7.5402e-14 as=3.0336e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.4338e-06 sim_w=5.76e-06 m_per_maxw=1.04167 numb_sub_cont=3 nfing=1 $X=310580 $Y=200 $D=22
M124 1 2 1 cpoly_n w=6e-06 l=2e-06 c=7.5402e-14 as=3.0336e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.4338e-06 sim_w=5.76e-06 m_per_maxw=1.04167 numb_sub_cont=3 nfing=1 $X=313100 $Y=200 $D=22
M125 1 2 1 cpoly_n w=6e-06 l=2e-06 c=7.5402e-14 as=3.0336e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.4338e-06 sim_w=5.76e-06 m_per_maxw=1.04167 numb_sub_cont=3 nfing=1 $X=315620 $Y=200 $D=22
M126 1 2 1 cpoly_n w=6e-06 l=2e-06 c=7.5402e-14 as=3.0336e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.4338e-06 sim_w=5.76e-06 m_per_maxw=1.04167 numb_sub_cont=3 nfing=1 $X=318140 $Y=200 $D=22
M127 1 2 1 cpoly_n w=6e-06 l=2e-06 c=7.5402e-14 as=3.0336e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.4338e-06 sim_w=5.76e-06 m_per_maxw=1.04167 numb_sub_cont=3 nfing=1 $X=320660 $Y=200 $D=22
M128 1 2 1 cpoly_n w=6e-06 l=2e-06 c=7.5402e-14 as=3.0336e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.4338e-06 sim_w=5.76e-06 m_per_maxw=1.04167 numb_sub_cont=3 nfing=1 $X=323180 $Y=200 $D=22
M129 1 2 1 cpoly_n w=6e-06 l=2e-06 c=7.5402e-14 as=3.0336e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.4338e-06 sim_w=5.76e-06 m_per_maxw=1.04167 numb_sub_cont=3 nfing=1 $X=325700 $Y=200 $D=22
M130 1 2 1 cpoly_n w=6e-06 l=2e-06 c=7.5402e-14 as=3.0336e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.4338e-06 sim_w=5.76e-06 m_per_maxw=1.04167 numb_sub_cont=3 nfing=1 $X=328220 $Y=200 $D=22
M131 1 2 1 cpoly_n w=6e-06 l=2e-06 c=7.5402e-14 as=3.0336e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.4338e-06 sim_w=5.76e-06 m_per_maxw=1.04167 numb_sub_cont=3 nfing=1 $X=330740 $Y=200 $D=22
M132 1 2 1 cpoly_n w=6e-06 l=2e-06 c=7.5402e-14 as=3.0336e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.4338e-06 sim_w=5.76e-06 m_per_maxw=1.04167 numb_sub_cont=3 nfing=1 $X=333260 $Y=200 $D=22
M133 1 2 1 cpoly_n w=6e-06 l=2e-06 c=7.5402e-14 as=3.0336e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.4338e-06 sim_w=5.76e-06 m_per_maxw=1.04167 numb_sub_cont=3 nfing=1 $X=335780 $Y=200 $D=22
M134 1 2 1 cpoly_n w=6e-06 l=2e-06 c=7.5402e-14 as=3.0336e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.4338e-06 sim_w=5.76e-06 m_per_maxw=1.04167 numb_sub_cont=3 nfing=1 $X=338300 $Y=200 $D=22
M135 1 2 1 cpoly_n w=6e-06 l=2e-06 c=7.5402e-14 as=3.0336e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.4338e-06 sim_w=5.76e-06 m_per_maxw=1.04167 numb_sub_cont=3 nfing=1 $X=340820 $Y=200 $D=22
M136 1 2 1 cpoly_n w=6e-06 l=2e-06 c=7.5402e-14 as=3.0336e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.4338e-06 sim_w=5.76e-06 m_per_maxw=1.04167 numb_sub_cont=3 nfing=1 $X=343340 $Y=200 $D=22
M137 1 2 1 cpoly_n w=6e-06 l=2e-06 c=7.5402e-14 as=3.0336e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.4338e-06 sim_w=5.76e-06 m_per_maxw=1.04167 numb_sub_cont=3 nfing=1 $X=345860 $Y=200 $D=22
M138 1 2 1 cpoly_n w=6e-06 l=2e-06 c=7.5402e-14 as=3.0336e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.4338e-06 sim_w=5.76e-06 m_per_maxw=1.04167 numb_sub_cont=3 nfing=1 $X=348380 $Y=200 $D=22
M139 1 2 1 cpoly_n w=6e-06 l=2e-06 c=7.5402e-14 as=3.0336e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.4338e-06 sim_w=5.76e-06 m_per_maxw=1.04167 numb_sub_cont=3 nfing=1 $X=350900 $Y=200 $D=22
M140 1 2 1 cpoly_n w=6e-06 l=2e-06 c=7.5402e-14 as=3.0336e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.4338e-06 sim_w=5.76e-06 m_per_maxw=1.04167 numb_sub_cont=3 nfing=1 $X=353420 $Y=200 $D=22
M141 1 2 1 cpoly_n w=6e-06 l=2e-06 c=7.5402e-14 as=3.0336e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.4338e-06 sim_w=5.76e-06 m_per_maxw=1.04167 numb_sub_cont=3 nfing=1 $X=355940 $Y=200 $D=22
M142 1 2 1 cpoly_n w=6e-06 l=2e-06 c=7.5402e-14 as=3.0336e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.4338e-06 sim_w=5.76e-06 m_per_maxw=1.04167 numb_sub_cont=3 nfing=1 $X=358460 $Y=200 $D=22
M143 1 2 1 cpoly_n w=6e-06 l=2e-06 c=7.5402e-14 as=3.0336e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.4338e-06 sim_w=5.76e-06 m_per_maxw=1.04167 numb_sub_cont=3 nfing=1 $X=360980 $Y=200 $D=22
M144 1 2 1 cpoly_n w=6e-06 l=2e-06 c=7.5402e-14 as=3.0336e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.4338e-06 sim_w=5.76e-06 m_per_maxw=1.04167 numb_sub_cont=3 nfing=1 $X=363500 $Y=200 $D=22
M145 1 2 1 cpoly_n w=6e-06 l=2e-06 c=7.5402e-14 as=3.0336e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.4338e-06 sim_w=5.76e-06 m_per_maxw=1.04167 numb_sub_cont=3 nfing=1 $X=366020 $Y=200 $D=22
M146 1 2 1 cpoly_n w=6e-06 l=2e-06 c=7.5402e-14 as=3.0336e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.4338e-06 sim_w=5.76e-06 m_per_maxw=1.04167 numb_sub_cont=3 nfing=1 $X=368540 $Y=200 $D=22
M147 1 2 1 cpoly_n w=6e-06 l=2e-06 c=7.5402e-14 as=3.0336e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.4338e-06 sim_w=5.76e-06 m_per_maxw=1.04167 numb_sub_cont=3 nfing=1 $X=371060 $Y=200 $D=22
M148 1 2 1 cpoly_n w=6e-06 l=2e-06 c=7.5402e-14 as=3.0336e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.4338e-06 sim_w=5.76e-06 m_per_maxw=1.04167 numb_sub_cont=3 nfing=1 $X=373580 $Y=200 $D=22
M149 1 2 1 cpoly_n w=6e-06 l=2e-06 c=7.5402e-14 as=3.0336e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.4338e-06 sim_w=5.76e-06 m_per_maxw=1.04167 numb_sub_cont=3 nfing=1 $X=376100 $Y=200 $D=22
M150 1 2 1 cpoly_n w=6e-06 l=2e-06 c=7.5402e-14 as=3.0336e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.4338e-06 sim_w=5.76e-06 m_per_maxw=1.04167 numb_sub_cont=3 nfing=1 $X=378620 $Y=200 $D=22
M151 1 2 1 cpoly_n w=6e-06 l=2e-06 c=7.5402e-14 as=3.0336e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.4338e-06 sim_w=5.76e-06 m_per_maxw=1.04167 numb_sub_cont=3 nfing=1 $X=381140 $Y=200 $D=22
M152 1 2 1 cpoly_n w=6e-06 l=2e-06 c=7.5402e-14 as=3.0336e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.4338e-06 sim_w=5.76e-06 m_per_maxw=1.04167 numb_sub_cont=3 nfing=1 $X=383660 $Y=200 $D=22
M153 1 2 1 cpoly_n w=6e-06 l=2e-06 c=7.5402e-14 as=3.0336e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.4338e-06 sim_w=5.76e-06 m_per_maxw=1.04167 numb_sub_cont=3 nfing=1 $X=386180 $Y=200 $D=22
M154 1 2 1 cpoly_n w=6e-06 l=2e-06 c=7.5402e-14 as=3.0336e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.4338e-06 sim_w=5.76e-06 m_per_maxw=1.04167 numb_sub_cont=3 nfing=1 $X=388700 $Y=200 $D=22
M155 1 2 1 cpoly_n w=6e-06 l=2e-06 c=7.5402e-14 as=3.0336e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.4338e-06 sim_w=5.76e-06 m_per_maxw=1.04167 numb_sub_cont=3 nfing=1 $X=391220 $Y=200 $D=22
M156 1 2 1 cpoly_n w=6e-06 l=2e-06 c=7.5402e-14 as=3.0336e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.4338e-06 sim_w=5.76e-06 m_per_maxw=1.04167 numb_sub_cont=3 nfing=1 $X=393740 $Y=200 $D=22
M157 1 2 1 cpoly_n w=6e-06 l=2e-06 c=7.5402e-14 as=3.0336e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.4338e-06 sim_w=5.76e-06 m_per_maxw=1.04167 numb_sub_cont=3 nfing=1 $X=396260 $Y=200 $D=22
M158 1 2 1 cpoly_n w=6e-06 l=2e-06 c=7.5402e-14 as=3.0336e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.4338e-06 sim_w=5.76e-06 m_per_maxw=1.04167 numb_sub_cont=3 nfing=1 $X=398780 $Y=200 $D=22
M159 1 2 1 cpoly_n w=6e-06 l=2e-06 c=7.5402e-14 as=3.0336e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.4338e-06 sim_w=5.76e-06 m_per_maxw=1.04167 numb_sub_cont=3 nfing=1 $X=401300 $Y=200 $D=22
M160 1 2 1 cpoly_n w=6e-06 l=2e-06 c=7.5402e-14 as=3.0336e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.4338e-06 sim_w=5.76e-06 m_per_maxw=1.04167 numb_sub_cont=3 nfing=1 $X=403820 $Y=200 $D=22
M161 1 2 1 cpoly_n w=6e-06 l=2e-06 c=7.5402e-14 as=3.0336e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.4338e-06 sim_w=5.76e-06 m_per_maxw=1.04167 numb_sub_cont=3 nfing=1 $X=406340 $Y=200 $D=22
M162 1 2 1 cpoly_n w=6e-06 l=2e-06 c=7.5402e-14 as=3.0336e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.4338e-06 sim_w=5.76e-06 m_per_maxw=1.04167 numb_sub_cont=3 nfing=1 $X=408860 $Y=200 $D=22
M163 1 2 1 cpoly_n w=6e-06 l=2e-06 c=7.5402e-14 as=2.4e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.4338e-06 sim_w=5.76e-06 m_per_maxw=1.04167 numb_sub_cont=3 nfing=1 $X=411380 $Y=200 $D=22
.ENDS
***************************************
.SUBCKT PAD_Fill_160 GND_PAD VDD_PAD gnd! vdd!
** N=5 EP=4 IP=26 FDC=1928
X0 gnd! vdd! cpoly_p_CDNS_58870478665105 $T=520 420500 0 0 $X=520 $Y=420500
X1 vdd! gnd! cpoly_n_CDNS_58870478665104 $T=520 433340 0 0 $X=520 $Y=433340
X2 GND_PAD VDD_PAD cpoly_p_CDNS_5887047866536 $T=15020 220 0 90 $X=7020 $Y=220
X3 GND_PAD VDD_PAD cpoly_p_CDNS_5887047866536 $T=43080 220 0 90 $X=35080 $Y=220
X4 GND_PAD VDD_PAD cpoly_p_CDNS_5887047866536 $T=71140 220 0 90 $X=63140 $Y=220
X5 GND_PAD VDD_PAD cpoly_p_CDNS_5887047866536 $T=99200 220 0 90 $X=91200 $Y=220
X6 GND_PAD VDD_PAD cpoly_p_CDNS_5887047866536 $T=127260 220 0 90 $X=119260 $Y=220
X7 GND_PAD VDD_PAD cpoly_p_CDNS_5887047866536 $T=155320 220 0 90 $X=147320 $Y=220
X8 VDD_PAD GND_PAD cpoly_n_CDNS_5887047866529 $T=28800 0 0 90 $X=21300 $Y=0
X9 VDD_PAD GND_PAD cpoly_n_CDNS_5887047866529 $T=56860 0 0 90 $X=49360 $Y=0
X10 VDD_PAD GND_PAD cpoly_n_CDNS_5887047866529 $T=84920 0 0 90 $X=77420 $Y=0
X11 VDD_PAD GND_PAD cpoly_n_CDNS_5887047866529 $T=112980 0 0 90 $X=105480 $Y=0
X12 VDD_PAD GND_PAD cpoly_n_CDNS_5887047866529 $T=141040 0 0 90 $X=133540 $Y=0
.ENDS
***************************************
.SUBCKT ICV_6 1 2
** N=2 EP=2 IP=2 FDC=164
X0 1 2 cpoly_p_CDNS_5887047866536 $T=0 0 0 0 $X=0 $Y=0
.ENDS
***************************************
.SUBCKT ICV_7 1 2
** N=2 EP=2 IP=2 FDC=164
X0 1 2 cpoly_p_CDNS_5887047866536 $T=0 0 0 0 $X=0 $Y=0
.ENDS
***************************************
.SUBCKT ICV_8 1 2
** N=2 EP=2 IP=2 FDC=164
X0 1 2 cpoly_p_CDNS_5887047866536 $T=0 0 0 0 $X=0 $Y=0
.ENDS
***************************************
.SUBCKT ICV_9 1 2
** N=2 EP=2 IP=2 FDC=164
X0 1 2 cpoly_p_CDNS_5887047866536 $T=0 0 0 0 $X=0 $Y=0
.ENDS
***************************************
.SUBCKT ICV_10 1 2
** N=2 EP=2 IP=2 FDC=164
X0 1 2 cpoly_p_CDNS_5887047866536 $T=0 0 0 0 $X=0 $Y=0
.ENDS
***************************************
.SUBCKT ICV_11 1 2
** N=2 EP=2 IP=2 FDC=164
X0 1 2 cpoly_p_CDNS_5887047866536 $T=0 0 0 0 $X=0 $Y=0
.ENDS
***************************************
.SUBCKT ICV_12 1 2
** N=2 EP=2 IP=2 FDC=164
X0 1 2 cpoly_p_CDNS_5887047866536 $T=0 0 0 0 $X=0 $Y=0
.ENDS
***************************************
.SUBCKT ICV_13 1 2
** N=2 EP=2 IP=2 FDC=164
X0 2 1 cpoly_n_CDNS_5887047866529 $T=0 0 0 0 $X=0 $Y=0
.ENDS
***************************************
.SUBCKT ICV_14 1 2
** N=2 EP=2 IP=2 FDC=164
X0 2 1 cpoly_n_CDNS_5887047866529 $T=0 0 0 0 $X=0 $Y=0
.ENDS
***************************************
.SUBCKT ICV_15 1 2
** N=2 EP=2 IP=2 FDC=164
X0 2 1 cpoly_n_CDNS_5887047866529 $T=0 0 0 0 $X=0 $Y=0
.ENDS
***************************************
.SUBCKT ICV_16 1 2
** N=2 EP=2 IP=2 FDC=164
X0 2 1 cpoly_n_CDNS_5887047866529 $T=0 0 0 0 $X=0 $Y=0
.ENDS
***************************************
.SUBCKT ICV_17 1 2
** N=2 EP=2 IP=2 FDC=164
X0 2 1 cpoly_n_CDNS_5887047866529 $T=0 0 0 0 $X=0 $Y=0
.ENDS
***************************************
.SUBCKT ICV_18 1 2
** N=2 EP=2 IP=2 FDC=164
X0 2 1 cpoly_n_CDNS_5887047866529 $T=0 0 0 0 $X=0 $Y=0
.ENDS
***************************************
.SUBCKT ICV_19 1 2
** N=2 EP=2 IP=2 FDC=164
X0 2 1 cpoly_n_CDNS_5887047866529 $T=0 0 0 0 $X=0 $Y=0
.ENDS
***************************************
.SUBCKT cpoly_p_CDNS_5887047866533 1 2
** N=2 EP=2 IP=0 FDC=78
M0 1 2 1 cpoly_p w=8.62e-06 l=2e-06 c=1.08536e-13 as=1.21314e-13 ad=7.488e-13 ps=1.44e-06 pd=1.21456e-06 sim_w=2.88e-06 m_per_maxw=2.99306 numb_sub_cont=4 nfing=1 $X=620 $Y=200 $D=21
M1 1 2 1 cpoly_p w=8.62e-06 l=2e-06 c=1.08536e-13 as=1.53388e-13 ad=7.488e-13 ps=1.44e-06 pd=1.21456e-06 sim_w=2.88e-06 m_per_maxw=2.99306 numb_sub_cont=4 nfing=1 $X=3140 $Y=200 $D=21
M2 1 2 1 cpoly_p w=8.62e-06 l=2e-06 c=1.08536e-13 as=1.53388e-13 ad=7.488e-13 ps=1.44e-06 pd=1.21456e-06 sim_w=2.88e-06 m_per_maxw=2.99306 numb_sub_cont=4 nfing=1 $X=5660 $Y=200 $D=21
M3 1 2 1 cpoly_p w=8.62e-06 l=2e-06 c=1.08536e-13 as=1.53388e-13 ad=7.488e-13 ps=1.44e-06 pd=1.21456e-06 sim_w=2.88e-06 m_per_maxw=2.99306 numb_sub_cont=4 nfing=1 $X=8180 $Y=200 $D=21
M4 1 2 1 cpoly_p w=8.62e-06 l=2e-06 c=1.08536e-13 as=1.53388e-13 ad=7.488e-13 ps=1.44e-06 pd=1.21456e-06 sim_w=2.88e-06 m_per_maxw=2.99306 numb_sub_cont=4 nfing=1 $X=10700 $Y=200 $D=21
M5 1 2 1 cpoly_p w=8.62e-06 l=2e-06 c=1.08536e-13 as=1.53388e-13 ad=7.488e-13 ps=1.44e-06 pd=1.21456e-06 sim_w=2.88e-06 m_per_maxw=2.99306 numb_sub_cont=4 nfing=1 $X=13220 $Y=200 $D=21
M6 1 2 1 cpoly_p w=8.62e-06 l=2e-06 c=1.08536e-13 as=1.53388e-13 ad=7.488e-13 ps=1.44e-06 pd=1.21456e-06 sim_w=2.88e-06 m_per_maxw=2.99306 numb_sub_cont=4 nfing=1 $X=15740 $Y=200 $D=21
M7 1 2 1 cpoly_p w=8.62e-06 l=2e-06 c=1.08536e-13 as=1.53388e-13 ad=7.488e-13 ps=1.44e-06 pd=1.21456e-06 sim_w=2.88e-06 m_per_maxw=2.99306 numb_sub_cont=4 nfing=1 $X=18260 $Y=200 $D=21
M8 1 2 1 cpoly_p w=8.62e-06 l=2e-06 c=1.08536e-13 as=1.53388e-13 ad=7.488e-13 ps=1.44e-06 pd=1.21456e-06 sim_w=2.88e-06 m_per_maxw=2.99306 numb_sub_cont=4 nfing=1 $X=20780 $Y=200 $D=21
M9 1 2 1 cpoly_p w=8.62e-06 l=2e-06 c=1.08536e-13 as=1.53388e-13 ad=7.488e-13 ps=1.44e-06 pd=1.21456e-06 sim_w=2.88e-06 m_per_maxw=2.99306 numb_sub_cont=4 nfing=1 $X=23300 $Y=200 $D=21
M10 1 2 1 cpoly_p w=8.62e-06 l=2e-06 c=1.08536e-13 as=1.53388e-13 ad=7.488e-13 ps=1.44e-06 pd=1.21456e-06 sim_w=2.88e-06 m_per_maxw=2.99306 numb_sub_cont=4 nfing=1 $X=25820 $Y=200 $D=21
M11 1 2 1 cpoly_p w=8.62e-06 l=2e-06 c=1.08536e-13 as=1.53388e-13 ad=7.488e-13 ps=1.44e-06 pd=1.21456e-06 sim_w=2.88e-06 m_per_maxw=2.99306 numb_sub_cont=4 nfing=1 $X=28340 $Y=200 $D=21
M12 1 2 1 cpoly_p w=8.62e-06 l=2e-06 c=1.08536e-13 as=1.53388e-13 ad=7.488e-13 ps=1.44e-06 pd=1.21456e-06 sim_w=2.88e-06 m_per_maxw=2.99306 numb_sub_cont=4 nfing=1 $X=30860 $Y=200 $D=21
M13 1 2 1 cpoly_p w=8.62e-06 l=2e-06 c=1.08536e-13 as=1.53388e-13 ad=7.488e-13 ps=1.44e-06 pd=1.21456e-06 sim_w=2.88e-06 m_per_maxw=2.99306 numb_sub_cont=4 nfing=1 $X=33380 $Y=200 $D=21
M14 1 2 1 cpoly_p w=8.62e-06 l=2e-06 c=1.08536e-13 as=1.53388e-13 ad=7.488e-13 ps=1.44e-06 pd=1.21456e-06 sim_w=2.88e-06 m_per_maxw=2.99306 numb_sub_cont=4 nfing=1 $X=35900 $Y=200 $D=21
M15 1 2 1 cpoly_p w=8.62e-06 l=2e-06 c=1.08536e-13 as=1.53388e-13 ad=7.488e-13 ps=1.44e-06 pd=1.21456e-06 sim_w=2.88e-06 m_per_maxw=2.99306 numb_sub_cont=4 nfing=1 $X=38420 $Y=200 $D=21
M16 1 2 1 cpoly_p w=8.62e-06 l=2e-06 c=1.08536e-13 as=1.53388e-13 ad=7.488e-13 ps=1.44e-06 pd=1.21456e-06 sim_w=2.88e-06 m_per_maxw=2.99306 numb_sub_cont=4 nfing=1 $X=40940 $Y=200 $D=21
M17 1 2 1 cpoly_p w=8.62e-06 l=2e-06 c=1.08536e-13 as=1.53388e-13 ad=7.488e-13 ps=1.44e-06 pd=1.21456e-06 sim_w=2.88e-06 m_per_maxw=2.99306 numb_sub_cont=4 nfing=1 $X=43460 $Y=200 $D=21
M18 1 2 1 cpoly_p w=8.62e-06 l=2e-06 c=1.08536e-13 as=1.53388e-13 ad=7.488e-13 ps=1.44e-06 pd=1.21456e-06 sim_w=2.88e-06 m_per_maxw=2.99306 numb_sub_cont=4 nfing=1 $X=45980 $Y=200 $D=21
M19 1 2 1 cpoly_p w=8.62e-06 l=2e-06 c=1.08536e-13 as=1.53388e-13 ad=7.488e-13 ps=1.44e-06 pd=1.21456e-06 sim_w=2.88e-06 m_per_maxw=2.99306 numb_sub_cont=4 nfing=1 $X=48500 $Y=200 $D=21
M20 1 2 1 cpoly_p w=8.62e-06 l=2e-06 c=1.08536e-13 as=1.53388e-13 ad=7.488e-13 ps=1.44e-06 pd=1.21456e-06 sim_w=2.88e-06 m_per_maxw=2.99306 numb_sub_cont=4 nfing=1 $X=51020 $Y=200 $D=21
M21 1 2 1 cpoly_p w=8.62e-06 l=2e-06 c=1.08536e-13 as=1.53388e-13 ad=7.488e-13 ps=1.44e-06 pd=1.21456e-06 sim_w=2.88e-06 m_per_maxw=2.99306 numb_sub_cont=4 nfing=1 $X=53540 $Y=200 $D=21
M22 1 2 1 cpoly_p w=8.62e-06 l=2e-06 c=1.08536e-13 as=1.53388e-13 ad=7.488e-13 ps=1.44e-06 pd=1.21456e-06 sim_w=2.88e-06 m_per_maxw=2.99306 numb_sub_cont=4 nfing=1 $X=56060 $Y=200 $D=21
M23 1 2 1 cpoly_p w=8.62e-06 l=2e-06 c=1.08536e-13 as=1.53388e-13 ad=7.488e-13 ps=1.44e-06 pd=1.21456e-06 sim_w=2.88e-06 m_per_maxw=2.99306 numb_sub_cont=4 nfing=1 $X=58580 $Y=200 $D=21
M24 1 2 1 cpoly_p w=8.62e-06 l=2e-06 c=1.08536e-13 as=1.53388e-13 ad=7.488e-13 ps=1.44e-06 pd=1.21456e-06 sim_w=2.88e-06 m_per_maxw=2.99306 numb_sub_cont=4 nfing=1 $X=61100 $Y=200 $D=21
M25 1 2 1 cpoly_p w=8.62e-06 l=2e-06 c=1.08536e-13 as=1.53388e-13 ad=7.488e-13 ps=1.44e-06 pd=1.21456e-06 sim_w=2.88e-06 m_per_maxw=2.99306 numb_sub_cont=4 nfing=1 $X=63620 $Y=200 $D=21
M26 1 2 1 cpoly_p w=8.62e-06 l=2e-06 c=1.08536e-13 as=1.53388e-13 ad=7.488e-13 ps=1.44e-06 pd=1.21456e-06 sim_w=2.88e-06 m_per_maxw=2.99306 numb_sub_cont=4 nfing=1 $X=66140 $Y=200 $D=21
M27 1 2 1 cpoly_p w=8.62e-06 l=2e-06 c=1.08536e-13 as=1.53388e-13 ad=7.488e-13 ps=1.44e-06 pd=1.21456e-06 sim_w=2.88e-06 m_per_maxw=2.99306 numb_sub_cont=4 nfing=1 $X=68660 $Y=200 $D=21
M28 1 2 1 cpoly_p w=8.62e-06 l=2e-06 c=1.08536e-13 as=1.53388e-13 ad=7.488e-13 ps=1.44e-06 pd=1.21456e-06 sim_w=2.88e-06 m_per_maxw=2.99306 numb_sub_cont=4 nfing=1 $X=71180 $Y=200 $D=21
M29 1 2 1 cpoly_p w=8.62e-06 l=2e-06 c=1.08536e-13 as=1.53388e-13 ad=7.488e-13 ps=1.44e-06 pd=1.21456e-06 sim_w=2.88e-06 m_per_maxw=2.99306 numb_sub_cont=4 nfing=1 $X=73700 $Y=200 $D=21
M30 1 2 1 cpoly_p w=8.62e-06 l=2e-06 c=1.08536e-13 as=1.53388e-13 ad=7.488e-13 ps=1.44e-06 pd=1.21456e-06 sim_w=2.88e-06 m_per_maxw=2.99306 numb_sub_cont=4 nfing=1 $X=76220 $Y=200 $D=21
M31 1 2 1 cpoly_p w=8.62e-06 l=2e-06 c=1.08536e-13 as=1.53388e-13 ad=7.488e-13 ps=1.44e-06 pd=1.21456e-06 sim_w=2.88e-06 m_per_maxw=2.99306 numb_sub_cont=4 nfing=1 $X=78740 $Y=200 $D=21
M32 1 2 1 cpoly_p w=8.62e-06 l=2e-06 c=1.08536e-13 as=1.53388e-13 ad=7.488e-13 ps=1.44e-06 pd=1.21456e-06 sim_w=2.88e-06 m_per_maxw=2.99306 numb_sub_cont=4 nfing=1 $X=81260 $Y=200 $D=21
M33 1 2 1 cpoly_p w=8.62e-06 l=2e-06 c=1.08536e-13 as=1.53388e-13 ad=7.488e-13 ps=1.44e-06 pd=1.21456e-06 sim_w=2.88e-06 m_per_maxw=2.99306 numb_sub_cont=4 nfing=1 $X=83780 $Y=200 $D=21
M34 1 2 1 cpoly_p w=8.62e-06 l=2e-06 c=1.08536e-13 as=1.53388e-13 ad=7.488e-13 ps=1.44e-06 pd=1.21456e-06 sim_w=2.88e-06 m_per_maxw=2.99306 numb_sub_cont=4 nfing=1 $X=86300 $Y=200 $D=21
M35 1 2 1 cpoly_p w=8.62e-06 l=2e-06 c=1.08536e-13 as=1.53388e-13 ad=7.488e-13 ps=1.44e-06 pd=1.21456e-06 sim_w=2.88e-06 m_per_maxw=2.99306 numb_sub_cont=4 nfing=1 $X=88820 $Y=200 $D=21
M36 1 2 1 cpoly_p w=8.62e-06 l=2e-06 c=1.08536e-13 as=1.53388e-13 ad=7.488e-13 ps=1.44e-06 pd=1.21456e-06 sim_w=2.88e-06 m_per_maxw=2.99306 numb_sub_cont=4 nfing=1 $X=91340 $Y=200 $D=21
M37 1 2 1 cpoly_p w=8.62e-06 l=2e-06 c=1.08536e-13 as=1.53388e-13 ad=7.488e-13 ps=1.44e-06 pd=1.21456e-06 sim_w=2.88e-06 m_per_maxw=2.99306 numb_sub_cont=4 nfing=1 $X=93860 $Y=200 $D=21
M38 1 2 1 cpoly_p w=8.62e-06 l=2e-06 c=1.08536e-13 as=1.53388e-13 ad=7.488e-13 ps=1.44e-06 pd=1.21456e-06 sim_w=2.88e-06 m_per_maxw=2.99306 numb_sub_cont=4 nfing=1 $X=96380 $Y=200 $D=21
M39 1 2 1 cpoly_p w=8.62e-06 l=2e-06 c=1.08536e-13 as=1.53388e-13 ad=7.488e-13 ps=1.44e-06 pd=1.21456e-06 sim_w=2.88e-06 m_per_maxw=2.99306 numb_sub_cont=4 nfing=1 $X=98900 $Y=200 $D=21
M40 1 2 1 cpoly_p w=8.62e-06 l=2e-06 c=1.08536e-13 as=1.53388e-13 ad=7.488e-13 ps=1.44e-06 pd=1.21456e-06 sim_w=2.88e-06 m_per_maxw=2.99306 numb_sub_cont=4 nfing=1 $X=101420 $Y=200 $D=21
M41 1 2 1 cpoly_p w=8.62e-06 l=2e-06 c=1.08536e-13 as=1.53388e-13 ad=7.488e-13 ps=1.44e-06 pd=1.21456e-06 sim_w=2.88e-06 m_per_maxw=2.99306 numb_sub_cont=4 nfing=1 $X=103940 $Y=200 $D=21
M42 1 2 1 cpoly_p w=8.62e-06 l=2e-06 c=1.08536e-13 as=1.53388e-13 ad=7.488e-13 ps=1.44e-06 pd=1.21456e-06 sim_w=2.88e-06 m_per_maxw=2.99306 numb_sub_cont=4 nfing=1 $X=106460 $Y=200 $D=21
M43 1 2 1 cpoly_p w=8.62e-06 l=2e-06 c=1.08536e-13 as=1.53388e-13 ad=7.488e-13 ps=1.44e-06 pd=1.21456e-06 sim_w=2.88e-06 m_per_maxw=2.99306 numb_sub_cont=4 nfing=1 $X=108980 $Y=200 $D=21
M44 1 2 1 cpoly_p w=8.62e-06 l=2e-06 c=1.08536e-13 as=1.53388e-13 ad=7.488e-13 ps=1.44e-06 pd=1.21456e-06 sim_w=2.88e-06 m_per_maxw=2.99306 numb_sub_cont=4 nfing=1 $X=111500 $Y=200 $D=21
M45 1 2 1 cpoly_p w=8.62e-06 l=2e-06 c=1.08536e-13 as=1.53388e-13 ad=7.488e-13 ps=1.44e-06 pd=1.21456e-06 sim_w=2.88e-06 m_per_maxw=2.99306 numb_sub_cont=4 nfing=1 $X=114020 $Y=200 $D=21
M46 1 2 1 cpoly_p w=8.62e-06 l=2e-06 c=1.08536e-13 as=1.53388e-13 ad=7.488e-13 ps=1.44e-06 pd=1.21456e-06 sim_w=2.88e-06 m_per_maxw=2.99306 numb_sub_cont=4 nfing=1 $X=116540 $Y=200 $D=21
M47 1 2 1 cpoly_p w=8.62e-06 l=2e-06 c=1.08536e-13 as=1.53388e-13 ad=7.488e-13 ps=1.44e-06 pd=1.21456e-06 sim_w=2.88e-06 m_per_maxw=2.99306 numb_sub_cont=4 nfing=1 $X=119060 $Y=200 $D=21
M48 1 2 1 cpoly_p w=8.62e-06 l=2e-06 c=1.08536e-13 as=1.53388e-13 ad=7.488e-13 ps=1.44e-06 pd=1.21456e-06 sim_w=2.88e-06 m_per_maxw=2.99306 numb_sub_cont=4 nfing=1 $X=121580 $Y=200 $D=21
M49 1 2 1 cpoly_p w=8.62e-06 l=2e-06 c=1.08536e-13 as=1.53388e-13 ad=7.488e-13 ps=1.44e-06 pd=1.21456e-06 sim_w=2.88e-06 m_per_maxw=2.99306 numb_sub_cont=4 nfing=1 $X=124100 $Y=200 $D=21
M50 1 2 1 cpoly_p w=8.62e-06 l=2e-06 c=1.08536e-13 as=1.53388e-13 ad=7.488e-13 ps=1.44e-06 pd=1.21456e-06 sim_w=2.88e-06 m_per_maxw=2.99306 numb_sub_cont=4 nfing=1 $X=126620 $Y=200 $D=21
M51 1 2 1 cpoly_p w=8.62e-06 l=2e-06 c=1.08536e-13 as=1.53388e-13 ad=7.488e-13 ps=1.44e-06 pd=1.21456e-06 sim_w=2.88e-06 m_per_maxw=2.99306 numb_sub_cont=4 nfing=1 $X=129140 $Y=200 $D=21
M52 1 2 1 cpoly_p w=8.62e-06 l=2e-06 c=1.08536e-13 as=1.53388e-13 ad=7.488e-13 ps=1.44e-06 pd=1.21456e-06 sim_w=2.88e-06 m_per_maxw=2.99306 numb_sub_cont=4 nfing=1 $X=131660 $Y=200 $D=21
M53 1 2 1 cpoly_p w=8.62e-06 l=2e-06 c=1.08536e-13 as=1.53388e-13 ad=7.488e-13 ps=1.44e-06 pd=1.21456e-06 sim_w=2.88e-06 m_per_maxw=2.99306 numb_sub_cont=4 nfing=1 $X=134180 $Y=200 $D=21
M54 1 2 1 cpoly_p w=8.62e-06 l=2e-06 c=1.08536e-13 as=1.53388e-13 ad=7.488e-13 ps=1.44e-06 pd=1.21456e-06 sim_w=2.88e-06 m_per_maxw=2.99306 numb_sub_cont=4 nfing=1 $X=136700 $Y=200 $D=21
M55 1 2 1 cpoly_p w=8.62e-06 l=2e-06 c=1.08536e-13 as=1.53388e-13 ad=7.488e-13 ps=1.44e-06 pd=1.21456e-06 sim_w=2.88e-06 m_per_maxw=2.99306 numb_sub_cont=4 nfing=1 $X=139220 $Y=200 $D=21
M56 1 2 1 cpoly_p w=8.62e-06 l=2e-06 c=1.08536e-13 as=1.53388e-13 ad=7.488e-13 ps=1.44e-06 pd=1.21456e-06 sim_w=2.88e-06 m_per_maxw=2.99306 numb_sub_cont=4 nfing=1 $X=141740 $Y=200 $D=21
M57 1 2 1 cpoly_p w=8.62e-06 l=2e-06 c=1.08536e-13 as=1.53388e-13 ad=7.488e-13 ps=1.44e-06 pd=1.21456e-06 sim_w=2.88e-06 m_per_maxw=2.99306 numb_sub_cont=4 nfing=1 $X=144260 $Y=200 $D=21
M58 1 2 1 cpoly_p w=8.62e-06 l=2e-06 c=1.08536e-13 as=1.53388e-13 ad=7.488e-13 ps=1.44e-06 pd=1.21456e-06 sim_w=2.88e-06 m_per_maxw=2.99306 numb_sub_cont=4 nfing=1 $X=146780 $Y=200 $D=21
M59 1 2 1 cpoly_p w=8.62e-06 l=2e-06 c=1.08536e-13 as=1.53388e-13 ad=7.488e-13 ps=1.44e-06 pd=1.21456e-06 sim_w=2.88e-06 m_per_maxw=2.99306 numb_sub_cont=4 nfing=1 $X=149300 $Y=200 $D=21
M60 1 2 1 cpoly_p w=8.62e-06 l=2e-06 c=1.08536e-13 as=1.53388e-13 ad=7.488e-13 ps=1.44e-06 pd=1.21456e-06 sim_w=2.88e-06 m_per_maxw=2.99306 numb_sub_cont=4 nfing=1 $X=151820 $Y=200 $D=21
M61 1 2 1 cpoly_p w=8.62e-06 l=2e-06 c=1.08536e-13 as=1.53388e-13 ad=7.488e-13 ps=1.44e-06 pd=1.21456e-06 sim_w=2.88e-06 m_per_maxw=2.99306 numb_sub_cont=4 nfing=1 $X=154340 $Y=200 $D=21
M62 1 2 1 cpoly_p w=8.62e-06 l=2e-06 c=1.08536e-13 as=1.53388e-13 ad=7.488e-13 ps=1.44e-06 pd=1.21456e-06 sim_w=2.88e-06 m_per_maxw=2.99306 numb_sub_cont=4 nfing=1 $X=156860 $Y=200 $D=21
M63 1 2 1 cpoly_p w=8.62e-06 l=2e-06 c=1.08536e-13 as=1.53388e-13 ad=7.488e-13 ps=1.44e-06 pd=1.21456e-06 sim_w=2.88e-06 m_per_maxw=2.99306 numb_sub_cont=4 nfing=1 $X=159380 $Y=200 $D=21
M64 1 2 1 cpoly_p w=8.62e-06 l=2e-06 c=1.08536e-13 as=1.53388e-13 ad=7.488e-13 ps=1.44e-06 pd=1.21456e-06 sim_w=2.88e-06 m_per_maxw=2.99306 numb_sub_cont=4 nfing=1 $X=161900 $Y=200 $D=21
M65 1 2 1 cpoly_p w=8.62e-06 l=2e-06 c=1.08536e-13 as=1.53388e-13 ad=7.488e-13 ps=1.44e-06 pd=1.21456e-06 sim_w=2.88e-06 m_per_maxw=2.99306 numb_sub_cont=4 nfing=1 $X=164420 $Y=200 $D=21
M66 1 2 1 cpoly_p w=8.62e-06 l=2e-06 c=1.08536e-13 as=1.53388e-13 ad=7.488e-13 ps=1.44e-06 pd=1.21456e-06 sim_w=2.88e-06 m_per_maxw=2.99306 numb_sub_cont=4 nfing=1 $X=166940 $Y=200 $D=21
M67 1 2 1 cpoly_p w=8.62e-06 l=2e-06 c=1.08536e-13 as=1.53388e-13 ad=7.488e-13 ps=1.44e-06 pd=1.21456e-06 sim_w=2.88e-06 m_per_maxw=2.99306 numb_sub_cont=4 nfing=1 $X=169460 $Y=200 $D=21
M68 1 2 1 cpoly_p w=8.62e-06 l=2e-06 c=1.08536e-13 as=1.53388e-13 ad=7.488e-13 ps=1.44e-06 pd=1.21456e-06 sim_w=2.88e-06 m_per_maxw=2.99306 numb_sub_cont=4 nfing=1 $X=171980 $Y=200 $D=21
M69 1 2 1 cpoly_p w=8.62e-06 l=2e-06 c=1.08536e-13 as=1.53388e-13 ad=7.488e-13 ps=1.44e-06 pd=1.21456e-06 sim_w=2.88e-06 m_per_maxw=2.99306 numb_sub_cont=4 nfing=1 $X=174500 $Y=200 $D=21
M70 1 2 1 cpoly_p w=8.62e-06 l=2e-06 c=1.08536e-13 as=1.53388e-13 ad=7.488e-13 ps=1.44e-06 pd=1.21456e-06 sim_w=2.88e-06 m_per_maxw=2.99306 numb_sub_cont=4 nfing=1 $X=177020 $Y=200 $D=21
M71 1 2 1 cpoly_p w=8.62e-06 l=2e-06 c=1.08536e-13 as=1.53388e-13 ad=7.488e-13 ps=1.44e-06 pd=1.21456e-06 sim_w=2.88e-06 m_per_maxw=2.99306 numb_sub_cont=4 nfing=1 $X=179540 $Y=200 $D=21
M72 1 2 1 cpoly_p w=8.62e-06 l=2e-06 c=1.08536e-13 as=1.53388e-13 ad=7.488e-13 ps=1.44e-06 pd=1.21456e-06 sim_w=2.88e-06 m_per_maxw=2.99306 numb_sub_cont=4 nfing=1 $X=182060 $Y=200 $D=21
M73 1 2 1 cpoly_p w=8.62e-06 l=2e-06 c=1.08536e-13 as=1.53388e-13 ad=7.488e-13 ps=1.44e-06 pd=1.21456e-06 sim_w=2.88e-06 m_per_maxw=2.99306 numb_sub_cont=4 nfing=1 $X=184580 $Y=200 $D=21
M74 1 2 1 cpoly_p w=8.62e-06 l=2e-06 c=1.08536e-13 as=1.53388e-13 ad=7.488e-13 ps=1.44e-06 pd=1.21456e-06 sim_w=2.88e-06 m_per_maxw=2.99306 numb_sub_cont=4 nfing=1 $X=187100 $Y=200 $D=21
M75 1 2 1 cpoly_p w=8.62e-06 l=2e-06 c=1.08536e-13 as=1.53388e-13 ad=7.488e-13 ps=1.44e-06 pd=1.21456e-06 sim_w=2.88e-06 m_per_maxw=2.99306 numb_sub_cont=4 nfing=1 $X=189620 $Y=200 $D=21
M76 1 2 1 cpoly_p w=8.62e-06 l=2e-06 c=1.08536e-13 as=1.53388e-13 ad=7.488e-13 ps=1.44e-06 pd=1.21456e-06 sim_w=2.88e-06 m_per_maxw=2.99306 numb_sub_cont=4 nfing=1 $X=192140 $Y=200 $D=21
M77 1 2 1 cpoly_p w=8.62e-06 l=2e-06 c=1.08536e-13 as=1.21314e-13 ad=7.488e-13 ps=1.44e-06 pd=1.21456e-06 sim_w=2.88e-06 m_per_maxw=2.99306 numb_sub_cont=4 nfing=1 $X=194660 $Y=200 $D=21
.ENDS
***************************************
.SUBCKT cpoly_n_CDNS_5887047866527 1 2
** N=2 EP=2 IP=0 FDC=78
M0 1 2 1 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=1.67141e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=620 $Y=200 $D=22
M1 1 2 1 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=3140 $Y=200 $D=22
M2 1 2 1 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=5660 $Y=200 $D=22
M3 1 2 1 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=8180 $Y=200 $D=22
M4 1 2 1 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=10700 $Y=200 $D=22
M5 1 2 1 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=13220 $Y=200 $D=22
M6 1 2 1 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=15740 $Y=200 $D=22
M7 1 2 1 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=18260 $Y=200 $D=22
M8 1 2 1 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=20780 $Y=200 $D=22
M9 1 2 1 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=23300 $Y=200 $D=22
M10 1 2 1 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=25820 $Y=200 $D=22
M11 1 2 1 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=28340 $Y=200 $D=22
M12 1 2 1 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=30860 $Y=200 $D=22
M13 1 2 1 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=33380 $Y=200 $D=22
M14 1 2 1 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=35900 $Y=200 $D=22
M15 1 2 1 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=38420 $Y=200 $D=22
M16 1 2 1 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=40940 $Y=200 $D=22
M17 1 2 1 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=43460 $Y=200 $D=22
M18 1 2 1 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=45980 $Y=200 $D=22
M19 1 2 1 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=48500 $Y=200 $D=22
M20 1 2 1 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=51020 $Y=200 $D=22
M21 1 2 1 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=53540 $Y=200 $D=22
M22 1 2 1 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=56060 $Y=200 $D=22
M23 1 2 1 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=58580 $Y=200 $D=22
M24 1 2 1 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=61100 $Y=200 $D=22
M25 1 2 1 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=63620 $Y=200 $D=22
M26 1 2 1 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=66140 $Y=200 $D=22
M27 1 2 1 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=68660 $Y=200 $D=22
M28 1 2 1 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=71180 $Y=200 $D=22
M29 1 2 1 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=73700 $Y=200 $D=22
M30 1 2 1 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=76220 $Y=200 $D=22
M31 1 2 1 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=78740 $Y=200 $D=22
M32 1 2 1 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=81260 $Y=200 $D=22
M33 1 2 1 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=83780 $Y=200 $D=22
M34 1 2 1 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=86300 $Y=200 $D=22
M35 1 2 1 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=88820 $Y=200 $D=22
M36 1 2 1 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=91340 $Y=200 $D=22
M37 1 2 1 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=93860 $Y=200 $D=22
M38 1 2 1 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=96380 $Y=200 $D=22
M39 1 2 1 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=98900 $Y=200 $D=22
M40 1 2 1 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=101420 $Y=200 $D=22
M41 1 2 1 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=103940 $Y=200 $D=22
M42 1 2 1 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=106460 $Y=200 $D=22
M43 1 2 1 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=108980 $Y=200 $D=22
M44 1 2 1 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=111500 $Y=200 $D=22
M45 1 2 1 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=114020 $Y=200 $D=22
M46 1 2 1 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=116540 $Y=200 $D=22
M47 1 2 1 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=119060 $Y=200 $D=22
M48 1 2 1 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=121580 $Y=200 $D=22
M49 1 2 1 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=124100 $Y=200 $D=22
M50 1 2 1 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=126620 $Y=200 $D=22
M51 1 2 1 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=129140 $Y=200 $D=22
M52 1 2 1 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=131660 $Y=200 $D=22
M53 1 2 1 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=134180 $Y=200 $D=22
M54 1 2 1 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=136700 $Y=200 $D=22
M55 1 2 1 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=139220 $Y=200 $D=22
M56 1 2 1 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=141740 $Y=200 $D=22
M57 1 2 1 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=144260 $Y=200 $D=22
M58 1 2 1 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=146780 $Y=200 $D=22
M59 1 2 1 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=149300 $Y=200 $D=22
M60 1 2 1 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=151820 $Y=200 $D=22
M61 1 2 1 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=154340 $Y=200 $D=22
M62 1 2 1 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=156860 $Y=200 $D=22
M63 1 2 1 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=159380 $Y=200 $D=22
M64 1 2 1 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=161900 $Y=200 $D=22
M65 1 2 1 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=164420 $Y=200 $D=22
M66 1 2 1 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=166940 $Y=200 $D=22
M67 1 2 1 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=169460 $Y=200 $D=22
M68 1 2 1 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=171980 $Y=200 $D=22
M69 1 2 1 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=174500 $Y=200 $D=22
M70 1 2 1 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=177020 $Y=200 $D=22
M71 1 2 1 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=179540 $Y=200 $D=22
M72 1 2 1 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=182060 $Y=200 $D=22
M73 1 2 1 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=184580 $Y=200 $D=22
M74 1 2 1 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=187100 $Y=200 $D=22
M75 1 2 1 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=189620 $Y=200 $D=22
M76 1 2 1 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=192140 $Y=200 $D=22
M77 1 2 1 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=1.67141e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=194660 $Y=200 $D=22
.ENDS
***************************************
.SUBCKT ICV_20 2 3
** N=4 EP=2 IP=4 FDC=156
X0 2 3 cpoly_p_CDNS_5887047866533 $T=520 420500 0 0 $X=520 $Y=420500
X1 3 2 cpoly_n_CDNS_5887047866527 $T=520 433340 0 0 $X=520 $Y=433340
.ENDS
***************************************
.SUBCKT ICV_21
** N=2 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT ICV_22
** N=2 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT ICV_23
** N=2 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT ICV_24
** N=2 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT ICV_25
** N=2 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT ICV_26
** N=3 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT ICV_27
** N=1 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT PAD_Fill_200 GND_PAD VDD_PAD gnd! vdd!
** N=5 EP=4 IP=46 FDC=2452
X0 GND_PAD VDD_PAD ICV_6 $T=183380 220 0 90 $X=175380 $Y=220
X1 GND_PAD VDD_PAD ICV_7 $T=155320 220 0 90 $X=147320 $Y=220
X2 GND_PAD VDD_PAD ICV_8 $T=127260 220 0 90 $X=119260 $Y=220
X3 GND_PAD VDD_PAD ICV_9 $T=99200 220 0 90 $X=91200 $Y=220
X4 GND_PAD VDD_PAD ICV_10 $T=71140 220 0 90 $X=63140 $Y=220
X5 GND_PAD VDD_PAD ICV_11 $T=43080 220 0 90 $X=35080 $Y=220
X6 GND_PAD VDD_PAD ICV_12 $T=15020 220 0 90 $X=7020 $Y=220
X7 GND_PAD VDD_PAD ICV_13 $T=197160 0 0 90 $X=189660 $Y=0
X8 GND_PAD VDD_PAD ICV_14 $T=169100 0 0 90 $X=161600 $Y=0
X9 GND_PAD VDD_PAD ICV_15 $T=141040 0 0 90 $X=133540 $Y=0
X10 GND_PAD VDD_PAD ICV_16 $T=112980 0 0 90 $X=105480 $Y=0
X11 GND_PAD VDD_PAD ICV_17 $T=84920 0 0 90 $X=77420 $Y=0
X12 GND_PAD VDD_PAD ICV_18 $T=56860 0 0 90 $X=49360 $Y=0
X13 GND_PAD VDD_PAD ICV_19 $T=28800 0 0 90 $X=21300 $Y=0
X14 gnd! vdd! ICV_20 $T=0 0 0 0 $X=0 $Y=371500
.ENDS
***************************************
.SUBCKT nOE_32 Bit_32 gnd! nOE Out vdd!
** N=7 EP=5 IP=0 FDC=6
M0 Out Bit_32 6 6 nmos_a L=2.4e-07 W=8e-07 AD=5.6e-13 AS=3.2e-13 PD=1.4e-06 PS=7e-07 w_cont=6e-07 nfing=1 source_num=2 $X=1040 $Y=320 $D=1
M1 6 7 gnd! gnd! nmos_a L=2.4e-07 W=8e-07 AD=5.6e-13 AS=3.2e-13 PD=1.4e-06 PS=7e-07 w_cont=6e-07 nfing=1 source_num=2 $X=2480 $Y=320 $D=1
M2 7 nOE gnd! gnd! nmos_a L=2.4e-07 W=4.8e-07 AD=4.32e-13 AS=1.92e-13 PD=1.08e-06 PS=5.4e-07 w_cont=6e-07 nfing=1 source_num=2 $X=4100 $Y=640 $D=1
M3 Out Bit_32 vdd! vdd! pmos_a L=2.4e-07 W=1e-06 AD=6.4e-13 AS=1.25e-13 PD=1.6e-06 PS=8e-07 w_cont=6e-07 nfing=1 mmm=1 $X=1040 $Y=2600 $D=5
M4 Out 7 vdd! vdd! pmos_a L=2.4e-07 W=1e-06 AD=6.4e-13 AS=1.25e-13 PD=1.6e-06 PS=8e-07 w_cont=6e-07 nfing=1 mmm=1 $X=2480 $Y=2600 $D=5
M5 7 nOE vdd! vdd! pmos_a L=2.4e-07 W=1e-06 AD=6.4e-13 AS=1.25e-13 PD=1.6e-06 PS=8e-07 w_cont=6e-07 nfing=1 mmm=1 $X=4100 $Y=2600 $D=5
.ENDS
***************************************
.SUBCKT nmos_a_CDNS_5887047866577
** N=3 EP=0 IP=0 FDC=0
*.SEEDPROM
.ENDS
***************************************
.SUBCKT pmos_a_CDNS_5887047866574 1 2 3
** N=3 EP=3 IP=0 FDC=2
M0 2 3 1 1 pmos_a L=2.4e-07 W=4e-06 AD=1.196e-12 AS=1.4e-13 PD=2.3e-06 PS=2.3e-06 w_cont=6e-07 nfing=1 mmm=1 $X=620 $Y=200 $D=5
M1 2 3 1 1 pmos_a L=2.4e-07 W=4e-06 AD=1.196e-12 AS=1.4e-13 PD=2.3e-06 PS=2.3e-06 w_cont=6e-07 nfing=1 mmm=1 $X=1380 $Y=200 $D=5
.ENDS
***************************************
.SUBCKT pmos_h_CDNS_5887047866578 1 2 3 4
** N=4 EP=4 IP=0 FDC=1
M0 3 4 2 1 pmos_h L=2.4e-07 W=1.5e-06 AD=6e-13 AS=6e-13 PD=2.3e-06 PS=2.3e-06 m=1 $X=820 $Y=600 $D=6
.ENDS
***************************************
.SUBCKT nmos_h_CDNS_5887047866576 1 2 3 4
** N=4 EP=4 IP=0 FDC=1
M0 3 4 2 1 nmos_h L=2.4e-07 W=7.2e-07 AD=2.88e-13 AS=2.88e-13 PD=1.52e-06 PS=1.52e-06 m=1 $X=820 $Y=600 $D=2
.ENDS
***************************************
.SUBCKT nmos_a_CDNS_5887047866572 1 2 3 4
** N=4 EP=4 IP=0 FDC=3
M0 2 3 1 1 nmos_a L=2.4e-07 W=2.4e-06 AD=9.1e-13 AS=9.6e-13 PD=1.75e-06 PS=1.75e-06 w_cont=1.1e-06 nfing=1 source_num=2 $X=620 $Y=200 $D=1
M1 2 3 1 1 nmos_a L=2.4e-07 W=2.4e-06 AD=9.1e-13 AS=1.248e-12 PD=1.75e-06 PS=1.75e-06 w_cont=1.1e-06 nfing=1 source_num=2 $X=1380 $Y=200 $D=1
M2 3 4 1 1 nmos_a L=2.4e-07 W=2.4e-06 AD=1.4e-12 AS=1.248e-12 PD=3.5e-06 PS=1.75e-06 w_cont=1.1e-06 nfing=1 source_num=2 $X=2140 $Y=200 $D=1
.ENDS
***************************************
.SUBCKT pmos_a_CDNS_5887047866575 1 2 3 4
** N=4 EP=4 IP=0 FDC=3
M0 2 3 1 1 pmos_a L=2.4e-07 W=4e-06 AD=1.196e-12 AS=1.4e-13 PD=2.3e-06 PS=2.3e-06 w_cont=6e-07 nfing=1 mmm=1 $X=620 $Y=200 $D=5
M1 2 3 1 1 pmos_a L=2.4e-07 W=4e-06 AD=1.196e-12 AS=1.76e-13 PD=2.3e-06 PS=2.3e-06 w_cont=6e-07 nfing=1 mmm=1 $X=1380 $Y=200 $D=5
M2 3 4 1 1 pmos_a L=2.4e-07 W=4e-06 AD=1.84e-12 AS=1.76e-13 PD=4.6e-06 PS=2.3e-06 w_cont=6e-07 nfing=1 mmm=1 $X=2140 $Y=200 $D=5
.ENDS
***************************************
.SUBCKT pmos_a_CDNS_5887047866579
** N=3 EP=0 IP=0 FDC=0
*.SEEDPROM
.ENDS
***************************************
.SUBCKT nmos_a_CDNS_5887047866573 1 2 3
** N=3 EP=3 IP=0 FDC=2
M0 2 3 1 1 nmos_a L=2.4e-07 W=2.4e-06 AD=9.1e-13 AS=9.6e-13 PD=1.75e-06 PS=1.75e-06 w_cont=1.1e-06 nfing=1 source_num=2 $X=620 $Y=200 $D=1
M1 2 3 1 1 nmos_a L=2.4e-07 W=2.4e-06 AD=9.1e-13 AS=9.6e-13 PD=1.75e-06 PS=1.75e-06 w_cont=1.1e-06 nfing=1 source_num=2 $X=1380 $Y=200 $D=1
.ENDS
***************************************
.SUBCKT Select_Bit Bit16 Bit32 A19 A18 DI_In DI_Out DI_Bank DO_Out DO_Bank DO_In vdd! gnd! In18 In19 High In16 In8 nA19 nA18 Low
** N=42 EP=20 IP=123 FDC=69
M0 22 22 gnd! gnd! nmos_a L=2.4e-07 W=6e-07 AD=4.8e-13 AS=2.4e-13 PD=1.2e-06 PS=6e-07 w_cont=6e-07 nfing=1 source_num=2 $X=-7180 $Y=580 $D=1
M1 23 26 gnd! gnd! nmos_a L=2.4e-07 W=6e-07 AD=4.8e-13 AS=2.4e-13 PD=1.2e-06 PS=6e-07 w_cont=6e-07 nfing=1 source_num=2 $X=-5360 $Y=-2240 $D=1
M2 26 Bit32 gnd! gnd! nmos_a L=2.4e-07 W=6e-07 AD=4.8e-13 AS=3.12e-13 PD=1.2e-06 PS=6e-07 w_cont=6e-07 nfing=1 source_num=2 $X=-3780 $Y=-3860 $D=1
M3 24 In16 gnd! gnd! nmos_a L=2.4e-07 W=6e-07 AD=4.8e-13 AS=3.12e-13 PD=1.2e-06 PS=6e-07 w_cont=6e-07 nfing=1 source_num=2 $X=-3780 $Y=-3100 $D=1
M4 26 Bit16 24 24 nmos_a L=2.4e-07 W=6e-07 AD=4.8e-13 AS=2.4e-13 PD=1.2e-06 PS=6e-07 w_cont=6e-07 nfing=1 source_num=2 $X=-3780 $Y=-1620 $D=1
M5 26 In8 gnd! gnd! nmos_a L=2.4e-07 W=6e-07 AD=4.8e-13 AS=3.12e-13 PD=1.2e-06 PS=6e-07 w_cont=6e-07 nfing=1 source_num=2 $X=-3780 $Y=-220 $D=1
M6 27 23 gnd! gnd! nmos_a L=2.4e-07 W=6e-07 AD=4.8e-13 AS=3.12e-13 PD=1.2e-06 PS=6e-07 w_cont=6e-07 nfing=1 source_num=2 $X=-3780 $Y=540 $D=1
M7 31 Bit16 gnd! gnd! nmos_a L=2.4e-07 W=6e-07 AD=4.8e-13 AS=2.4e-13 PD=1.2e-06 PS=6e-07 w_cont=6e-07 nfing=1 source_num=2 $X=2840 $Y=-2020 $D=1
M8 31 Bit32 gnd! gnd! nmos_a L=2.4e-07 W=6e-07 AD=4.8e-13 AS=3.12e-13 PD=1.2e-06 PS=6e-07 w_cont=6e-07 nfing=1 source_num=2 $X=4320 $Y=-2020 $D=1
M9 32 31 gnd! gnd! nmos_a L=2.4e-07 W=6e-07 AD=4.8e-13 AS=3.12e-13 PD=1.2e-06 PS=6e-07 w_cont=6e-07 nfing=1 source_num=2 $X=5080 $Y=-2020 $D=1
M10 36 34 gnd! gnd! nmos_a L=2.4e-07 W=6e-07 AD=3.12e-13 AS=2.4e-13 PD=6e-07 PS=6e-07 w_cont=6e-07 nfing=1 source_num=2 $X=8840 $Y=-2020 $D=1
M11 36 In19 gnd! gnd! nmos_a L=2.4e-07 W=6e-07 AD=3.12e-13 AS=2.4e-13 PD=6e-07 PS=6e-07 w_cont=6e-07 nfing=1 source_num=2 $X=9600 $Y=-2020 $D=1
M12 40 36 gnd! gnd! nmos_a L=2.4e-07 W=6e-07 AD=4.8e-13 AS=3.12e-13 PD=1.2e-06 PS=6e-07 w_cont=6e-07 nfing=1 source_num=2 $X=11220 $Y=-2020 $D=1
M13 Low High gnd! gnd! nmos_a L=2.4e-07 W=6e-07 AD=4.8e-13 AS=2.4e-13 PD=1.2e-06 PS=6e-07 w_cont=6e-07 nfing=1 source_num=2 $X=-7480 $Y=-5340 $D=1
M14 34 In18 32 32 nmos_a L=2.4e-07 W=6e-07 AD=4.8e-13 AS=2.4e-13 PD=1.2e-06 PS=6e-07 w_cont=6e-07 nfing=1 source_num=2 $X=6520 $Y=-2020 $D=1
M15 37 40 gnd! gnd! nmos_a L=2.4e-07 W=6e-07 AD=4.8e-13 AS=2.4e-13 PD=1.2e-06 PS=6e-07 w_cont=6e-07 nfing=1 source_num=2 $X=10920 $Y=540 $D=1
M16 40 41 gnd! gnd! nmos_a L=2.4e-07 W=6e-07 AD=4.8e-13 AS=3.12e-13 PD=1.2e-06 PS=6e-07 w_cont=6e-07 nfing=1 source_num=2 $X=11980 $Y=-2020 $D=1
M17 41 In18 gnd! gnd! nmos_a L=2.4e-07 W=6e-07 AD=4.8e-13 AS=3.12e-13 PD=1.2e-06 PS=6e-07 w_cont=6e-07 nfing=1 source_num=2 $X=14080 $Y=-2020 $D=1
M18 41 Bit32 gnd! gnd! nmos_a L=2.4e-07 W=6e-07 AD=4.8e-13 AS=3.12e-13 PD=1.2e-06 PS=6e-07 w_cont=6e-07 nfing=1 source_num=2 $X=14840 $Y=-2020 $D=1
M19 nA19 A19 gnd! gnd! nmos_a L=2.4e-07 W=6e-07 AD=4.8e-13 AS=2.4e-13 PD=1.2e-06 PS=6e-07 w_cont=6e-07 nfing=1 source_num=2 $X=17000 $Y=-5400 $D=1
M20 nA18 A18 gnd! gnd! nmos_a L=2.4e-07 W=6e-07 AD=4.8e-13 AS=2.4e-13 PD=1.2e-06 PS=6e-07 w_cont=6e-07 nfing=1 source_num=2 $X=17000 $Y=3500 $D=1
M21 23 26 vdd! vdd! pmos_a L=2.4e-07 W=1.2e-06 AD=7.2e-13 AS=1.26e-13 PD=1.8e-06 PS=9e-07 w_cont=6e-07 nfing=1 mmm=1 $X=-5360 $Y=-4440 $D=5
M22 26 Bit32 28 28 pmos_a L=2.4e-07 W=1.2e-06 AD=7.2e-13 AS=1.26e-13 PD=1.8e-06 PS=9e-07 w_cont=6e-07 nfing=1 mmm=1 $X=-1880 $Y=-4540 $D=5
M23 28 In16 29 29 pmos_a L=2.4e-07 W=1.2e-06 AD=7.2e-13 AS=1.62e-13 PD=1.8e-06 PS=9e-07 w_cont=6e-07 nfing=1 mmm=1 $X=-1880 $Y=-3100 $D=5
M24 28 Bit16 29 29 pmos_a L=2.4e-07 W=1.2e-06 AD=7.2e-13 AS=1.62e-13 PD=1.8e-06 PS=9e-07 w_cont=6e-07 nfing=1 mmm=1 $X=-1880 $Y=-2340 $D=5
M25 29 In8 vdd! vdd! pmos_a L=2.4e-07 W=1.2e-06 AD=7.2e-13 AS=1.26e-13 PD=1.8e-06 PS=9e-07 w_cont=6e-07 nfing=1 mmm=1 $X=-1880 $Y=-940 $D=5
M26 27 23 vdd! vdd! pmos_a L=2.4e-07 W=1e-06 AD=6.4e-13 AS=1.25e-13 PD=1.6e-06 PS=8e-07 w_cont=6e-07 nfing=1 mmm=1 $X=-1680 $Y=540 $D=5
M27 36 In19 35 35 pmos_a L=2.4e-07 W=2e-06 AD=1.04e-12 AS=1.3e-13 PD=2.6e-06 PS=1.3e-06 w_cont=6e-07 nfing=1 mmm=1 $X=9600 $Y=-5400 $D=5
M28 30 Bit16 vdd! vdd! pmos_a L=2.4e-07 W=2e-06 AD=1.04e-12 AS=1.3e-13 PD=2.6e-06 PS=1.3e-06 w_cont=6e-07 nfing=1 mmm=1 $X=2840 $Y=-5020 $D=5
M29 31 Bit32 30 30 pmos_a L=2.4e-07 W=2e-06 AD=1.04e-12 AS=1.3e-13 PD=2.6e-06 PS=1.3e-06 w_cont=6e-07 nfing=1 mmm=1 $X=4320 $Y=-5400 $D=5
M30 35 34 vdd! vdd! pmos_a L=2.4e-07 W=2e-06 AD=1.04e-12 AS=1.3e-13 PD=2.6e-06 PS=1.3e-06 w_cont=6e-07 nfing=1 mmm=1 $X=8160 $Y=-5400 $D=5
M31 39 36 vdd! vdd! pmos_a L=2.4e-07 W=2e-06 AD=1.04e-12 AS=1.3e-13 PD=2.6e-06 PS=1.3e-06 w_cont=6e-07 nfing=1 mmm=1 $X=11040 $Y=-5400 $D=5
M32 40 41 39 39 pmos_a L=2.4e-07 W=2e-06 AD=1.04e-12 AS=1.3e-13 PD=2.6e-06 PS=1.3e-06 w_cont=6e-07 nfing=1 mmm=1 $X=12480 $Y=-5400 $D=5
M33 42 In18 vdd! vdd! pmos_a L=2.4e-07 W=2e-06 AD=1.04e-12 AS=1.3e-13 PD=2.6e-06 PS=1.3e-06 w_cont=6e-07 nfing=1 mmm=1 $X=13920 $Y=-5400 $D=5
M34 41 Bit32 42 42 pmos_a L=2.4e-07 W=2e-06 AD=1.04e-12 AS=1.3e-13 PD=2.6e-06 PS=1.3e-06 w_cont=6e-07 nfing=1 mmm=1 $X=15360 $Y=-5400 $D=5
M35 37 40 vdd! vdd! pmos_a L=2.4e-07 W=1e-06 AD=6.4e-13 AS=1.25e-13 PD=1.6e-06 PS=8e-07 w_cont=6e-07 nfing=1 mmm=1 $X=8360 $Y=540 $D=5
M36 High 22 vdd! vdd! pmos_a L=2.4e-07 W=6e-07 AD=4.8e-13 AS=1.23e-13 PD=1.2e-06 PS=6e-07 w_cont=6e-07 nfing=1 mmm=1 $X=-7480 $Y=-1840 $D=5
M37 34 31 vdd! vdd! pmos_a L=2.4e-07 W=6e-07 AD=4.8e-13 AS=1.59e-13 PD=1.2e-06 PS=6e-07 w_cont=6e-07 nfing=1 mmm=1 $X=5760 $Y=-4620 $D=5
M38 34 In18 vdd! vdd! pmos_a L=2.4e-07 W=6e-07 AD=4.8e-13 AS=1.59e-13 PD=1.2e-06 PS=6e-07 w_cont=6e-07 nfing=1 mmm=1 $X=6520 $Y=-4620 $D=5
X39 vdd! nA19 A19 pmos_a_CDNS_5887047866540 $T=17860 -1300 0 180 $X=16420 $Y=-3500
X40 vdd! nA18 A18 pmos_a_CDNS_5887047866540 $T=17860 7720 0 180 $X=16420 $Y=5520
X57 vdd! DI_Bank 25 pmos_a_CDNS_5887047866574 $T=-7700 4380 0 0 $X=-7700 $Y=4380
X58 vdd! DO_Out 38 pmos_a_CDNS_5887047866574 $T=15780 4380 1 180 $X=13540 $Y=4380
X59 vdd! DI_Out 21 23 pmos_h_CDNS_5887047866578 $T=-4920 1680 1 180 $X=-8060 $Y=1680
X60 vdd! DI_In 21 27 pmos_h_CDNS_5887047866578 $T=580 1680 1 180 $X=-2560 $Y=1680
X61 vdd! DO_Bank 33 37 pmos_h_CDNS_5887047866578 $T=7500 1680 0 0 $X=7500 $Y=1680
X62 vdd! DO_In 33 40 pmos_h_CDNS_5887047866578 $T=13000 1680 0 0 $X=13000 $Y=1680
X63 gnd! DI_Out 21 27 nmos_h_CDNS_5887047866576 $T=-2560 1680 1 180 $X=-4920 $Y=1680
X64 gnd! DI_In 21 23 nmos_h_CDNS_5887047866576 $T=2940 2060 1 180 $X=580 $Y=2060
X65 gnd! DO_Bank 33 40 nmos_h_CDNS_5887047866576 $T=5140 1680 0 0 $X=5140 $Y=1680
X66 gnd! DO_In 33 37 nmos_h_CDNS_5887047866576 $T=10640 1680 0 0 $X=10640 $Y=1680
X67 gnd! DI_Bank 25 21 nmos_a_CDNS_5887047866572 $T=-5460 4960 0 0 $X=-5460 $Y=4960
X68 gnd! DO_Out 38 33 nmos_a_CDNS_5887047866572 $T=13540 4960 1 180 $X=10580 $Y=4960
X69 vdd! DI_Bank 25 21 pmos_a_CDNS_5887047866575 $T=460 4380 1 180 $X=-2500 $Y=4380
X70 vdd! DO_Out 38 33 pmos_a_CDNS_5887047866575 $T=7620 4380 0 0 $X=7620 $Y=4380
X74 gnd! DI_Bank 25 nmos_a_CDNS_5887047866573 $T=460 4960 0 0 $X=460 $Y=4960
X75 gnd! DO_Out 38 nmos_a_CDNS_5887047866573 $T=7620 4960 1 180 $X=5380 $Y=4960
.ENDS
***************************************
.SUBCKT Cell1 gnd! vdd! nW High 12
** N=12 EP=5 IP=0 FDC=5
*.SEEDPROM
M0 High 12 gnd! gnd! nmos_a L=3.8e-07 W=4.8e-07 AD=9.258e-13 AS=2.496e-13 PD=1.06e-06 PS=5.3e-07 w_cont=5.8e-07 nfing=1 source_num=2 $X=260 $Y=3520 $D=1
M1 High 12 vdd! vdd! pmos_a L=2.4e-07 W=1e-06 AD=5.928e-13 AS=1.25e-13 PD=1.6e-06 PS=8e-07 w_cont=6e-07 nfing=1 mmm=1 $X=700 $Y=5300 $D=5
M2 12 High gnd! gnd! pmos_a L=2.4e-07 W=1e-06 AD=5.928e-13 AS=1.25e-13 PD=1.6e-06 PS=8e-07 w_cont=6e-07 nfing=1 mmm=1 $X=900 $Y=260 $D=5
M3 Data nW High vdd! pmos_h L=2.4e-07 W=6.6e-07 AD=2.64e-13 AS=2.64e-13 PD=1.46e-06 PS=1.46e-06 m=1 $X=600 $Y=1860 $D=6
M4 12 nW nData vdd! pmos_h L=2.4e-07 W=6.6e-07 AD=2.64e-13 AS=2.64e-13 PD=1.46e-06 PS=1.46e-06 m=1 $X=2360 $Y=3280 $D=6
.ENDS
***************************************
.SUBCKT ICV_28 4 5 7 8 9 10
** N=10 EP=6 IP=20 FDC=10
*.SEEDPROM
X0 4 5 5 7 8 Cell1 $T=0 0 1 180 $X=-3560 $Y=-440
X1 4 5 5 9 10 Cell1 $T=0 0 0 0 $X=-320 $Y=-440
.ENDS
***************************************
.SUBCKT ICV_29 4 5 7 8 9 10
** N=14 EP=6 IP=20 FDC=22
*.SEEDPROM
M0 12 11 4 4 nmos_a L=3.8e-07 W=4.8e-07 AD=9.258e-13 AS=2.496e-13 PD=1.06e-06 PS=5.3e-07 w_cont=5.8e-07 nfing=1 source_num=2 $X=-3840 $Y=1220 $D=1
M1 14 13 4 4 nmos_a L=3.8e-07 W=4.8e-07 AD=9.258e-13 AS=2.496e-13 PD=1.06e-06 PS=5.3e-07 w_cont=5.8e-07 nfing=1 source_num=2 $X=-2940 $Y=1220 $D=1
X2 4 5 7 8 11 12 ICV_28 $T=-6400 0 0 0 $X=-9960 $Y=-440
X3 4 5 13 14 9 10 ICV_28 $T=0 0 0 0 $X=-3560 $Y=-440
.ENDS
***************************************
.SUBCKT cpoly_p_CDNS_58870478665103 1 2
** N=2 EP=2 IP=0 FDC=20
M0 1 2 1 cpoly_p w=6e-06 l=2e-06 c=8.0712e-14 as=1.68e-13 ad=7.488e-13 ps=1.44e-06 pd=1.13684e-06 sim_w=2.88e-06 m_per_maxw=2.08333 numb_sub_cont=4 nfing=1 $X=620 $Y=200 $D=21
M1 1 2 1 cpoly_p w=6e-06 l=2e-06 c=8.0712e-14 as=2.1408e-13 ad=7.488e-13 ps=1.44e-06 pd=1.13684e-06 sim_w=2.88e-06 m_per_maxw=2.08333 numb_sub_cont=4 nfing=1 $X=3140 $Y=200 $D=21
M2 1 2 1 cpoly_p w=6e-06 l=2e-06 c=8.0712e-14 as=2.1408e-13 ad=7.488e-13 ps=1.44e-06 pd=1.13684e-06 sim_w=2.88e-06 m_per_maxw=2.08333 numb_sub_cont=4 nfing=1 $X=5660 $Y=200 $D=21
M3 1 2 1 cpoly_p w=6e-06 l=2e-06 c=8.0712e-14 as=2.1408e-13 ad=7.488e-13 ps=1.44e-06 pd=1.13684e-06 sim_w=2.88e-06 m_per_maxw=2.08333 numb_sub_cont=4 nfing=1 $X=8180 $Y=200 $D=21
M4 1 2 1 cpoly_p w=6e-06 l=2e-06 c=8.0712e-14 as=2.1408e-13 ad=7.488e-13 ps=1.44e-06 pd=1.13684e-06 sim_w=2.88e-06 m_per_maxw=2.08333 numb_sub_cont=4 nfing=1 $X=10700 $Y=200 $D=21
M5 1 2 1 cpoly_p w=6e-06 l=2e-06 c=8.0712e-14 as=2.1408e-13 ad=7.488e-13 ps=1.44e-06 pd=1.13684e-06 sim_w=2.88e-06 m_per_maxw=2.08333 numb_sub_cont=4 nfing=1 $X=13220 $Y=200 $D=21
M6 1 2 1 cpoly_p w=6e-06 l=2e-06 c=8.0712e-14 as=2.1408e-13 ad=7.488e-13 ps=1.44e-06 pd=1.13684e-06 sim_w=2.88e-06 m_per_maxw=2.08333 numb_sub_cont=4 nfing=1 $X=15740 $Y=200 $D=21
M7 1 2 1 cpoly_p w=6e-06 l=2e-06 c=8.0712e-14 as=2.1408e-13 ad=7.488e-13 ps=1.44e-06 pd=1.13684e-06 sim_w=2.88e-06 m_per_maxw=2.08333 numb_sub_cont=4 nfing=1 $X=18260 $Y=200 $D=21
M8 1 2 1 cpoly_p w=6e-06 l=2e-06 c=8.0712e-14 as=2.1408e-13 ad=7.488e-13 ps=1.44e-06 pd=1.13684e-06 sim_w=2.88e-06 m_per_maxw=2.08333 numb_sub_cont=4 nfing=1 $X=20780 $Y=200 $D=21
M9 1 2 1 cpoly_p w=6e-06 l=2e-06 c=8.0712e-14 as=2.1408e-13 ad=7.488e-13 ps=1.44e-06 pd=1.13684e-06 sim_w=2.88e-06 m_per_maxw=2.08333 numb_sub_cont=4 nfing=1 $X=23300 $Y=200 $D=21
M10 1 2 1 cpoly_p w=6e-06 l=2e-06 c=8.0712e-14 as=2.1408e-13 ad=7.488e-13 ps=1.44e-06 pd=1.13684e-06 sim_w=2.88e-06 m_per_maxw=2.08333 numb_sub_cont=4 nfing=1 $X=25820 $Y=200 $D=21
M11 1 2 1 cpoly_p w=6e-06 l=2e-06 c=8.0712e-14 as=2.1408e-13 ad=7.488e-13 ps=1.44e-06 pd=1.13684e-06 sim_w=2.88e-06 m_per_maxw=2.08333 numb_sub_cont=4 nfing=1 $X=28340 $Y=200 $D=21
M12 1 2 1 cpoly_p w=6e-06 l=2e-06 c=8.0712e-14 as=2.1408e-13 ad=7.488e-13 ps=1.44e-06 pd=1.13684e-06 sim_w=2.88e-06 m_per_maxw=2.08333 numb_sub_cont=4 nfing=1 $X=30860 $Y=200 $D=21
M13 1 2 1 cpoly_p w=6e-06 l=2e-06 c=8.0712e-14 as=2.1408e-13 ad=7.488e-13 ps=1.44e-06 pd=1.13684e-06 sim_w=2.88e-06 m_per_maxw=2.08333 numb_sub_cont=4 nfing=1 $X=33380 $Y=200 $D=21
M14 1 2 1 cpoly_p w=6e-06 l=2e-06 c=8.0712e-14 as=2.1408e-13 ad=7.488e-13 ps=1.44e-06 pd=1.13684e-06 sim_w=2.88e-06 m_per_maxw=2.08333 numb_sub_cont=4 nfing=1 $X=35900 $Y=200 $D=21
M15 1 2 1 cpoly_p w=6e-06 l=2e-06 c=8.0712e-14 as=2.1408e-13 ad=7.488e-13 ps=1.44e-06 pd=1.13684e-06 sim_w=2.88e-06 m_per_maxw=2.08333 numb_sub_cont=4 nfing=1 $X=38420 $Y=200 $D=21
M16 1 2 1 cpoly_p w=6e-06 l=2e-06 c=8.0712e-14 as=2.1408e-13 ad=7.488e-13 ps=1.44e-06 pd=1.13684e-06 sim_w=2.88e-06 m_per_maxw=2.08333 numb_sub_cont=4 nfing=1 $X=40940 $Y=200 $D=21
M17 1 2 1 cpoly_p w=6e-06 l=2e-06 c=8.0712e-14 as=2.1408e-13 ad=7.488e-13 ps=1.44e-06 pd=1.13684e-06 sim_w=2.88e-06 m_per_maxw=2.08333 numb_sub_cont=4 nfing=1 $X=43460 $Y=200 $D=21
M18 1 2 1 cpoly_p w=6e-06 l=2e-06 c=8.0712e-14 as=2.1408e-13 ad=7.488e-13 ps=1.44e-06 pd=1.13684e-06 sim_w=2.88e-06 m_per_maxw=2.08333 numb_sub_cont=4 nfing=1 $X=45980 $Y=200 $D=21
M19 1 2 1 cpoly_p w=6e-06 l=2e-06 c=8.0712e-14 as=1.68e-13 ad=7.488e-13 ps=1.44e-06 pd=1.13684e-06 sim_w=2.88e-06 m_per_maxw=2.08333 numb_sub_cont=4 nfing=1 $X=48500 $Y=200 $D=21
.ENDS
***************************************
.SUBCKT cpoly_n_CDNS_58870478665102 1 2
** N=2 EP=2 IP=0 FDC=20
M0 1 2 1 cpoly_n w=6e-06 l=2e-06 c=7.5402e-14 as=2.4e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.4338e-06 sim_w=5.76e-06 m_per_maxw=1.04167 numb_sub_cont=3 nfing=1 $X=620 $Y=200 $D=22
M1 1 2 1 cpoly_n w=6e-06 l=2e-06 c=7.5402e-14 as=3.0336e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.4338e-06 sim_w=5.76e-06 m_per_maxw=1.04167 numb_sub_cont=3 nfing=1 $X=3140 $Y=200 $D=22
M2 1 2 1 cpoly_n w=6e-06 l=2e-06 c=7.5402e-14 as=3.0336e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.4338e-06 sim_w=5.76e-06 m_per_maxw=1.04167 numb_sub_cont=3 nfing=1 $X=5660 $Y=200 $D=22
M3 1 2 1 cpoly_n w=6e-06 l=2e-06 c=7.5402e-14 as=3.0336e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.4338e-06 sim_w=5.76e-06 m_per_maxw=1.04167 numb_sub_cont=3 nfing=1 $X=8180 $Y=200 $D=22
M4 1 2 1 cpoly_n w=6e-06 l=2e-06 c=7.5402e-14 as=3.0336e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.4338e-06 sim_w=5.76e-06 m_per_maxw=1.04167 numb_sub_cont=3 nfing=1 $X=10700 $Y=200 $D=22
M5 1 2 1 cpoly_n w=6e-06 l=2e-06 c=7.5402e-14 as=3.0336e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.4338e-06 sim_w=5.76e-06 m_per_maxw=1.04167 numb_sub_cont=3 nfing=1 $X=13220 $Y=200 $D=22
M6 1 2 1 cpoly_n w=6e-06 l=2e-06 c=7.5402e-14 as=3.0336e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.4338e-06 sim_w=5.76e-06 m_per_maxw=1.04167 numb_sub_cont=3 nfing=1 $X=15740 $Y=200 $D=22
M7 1 2 1 cpoly_n w=6e-06 l=2e-06 c=7.5402e-14 as=3.0336e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.4338e-06 sim_w=5.76e-06 m_per_maxw=1.04167 numb_sub_cont=3 nfing=1 $X=18260 $Y=200 $D=22
M8 1 2 1 cpoly_n w=6e-06 l=2e-06 c=7.5402e-14 as=3.0336e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.4338e-06 sim_w=5.76e-06 m_per_maxw=1.04167 numb_sub_cont=3 nfing=1 $X=20780 $Y=200 $D=22
M9 1 2 1 cpoly_n w=6e-06 l=2e-06 c=7.5402e-14 as=3.0336e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.4338e-06 sim_w=5.76e-06 m_per_maxw=1.04167 numb_sub_cont=3 nfing=1 $X=23300 $Y=200 $D=22
M10 1 2 1 cpoly_n w=6e-06 l=2e-06 c=7.5402e-14 as=3.0336e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.4338e-06 sim_w=5.76e-06 m_per_maxw=1.04167 numb_sub_cont=3 nfing=1 $X=25820 $Y=200 $D=22
M11 1 2 1 cpoly_n w=6e-06 l=2e-06 c=7.5402e-14 as=3.0336e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.4338e-06 sim_w=5.76e-06 m_per_maxw=1.04167 numb_sub_cont=3 nfing=1 $X=28340 $Y=200 $D=22
M12 1 2 1 cpoly_n w=6e-06 l=2e-06 c=7.5402e-14 as=3.0336e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.4338e-06 sim_w=5.76e-06 m_per_maxw=1.04167 numb_sub_cont=3 nfing=1 $X=30860 $Y=200 $D=22
M13 1 2 1 cpoly_n w=6e-06 l=2e-06 c=7.5402e-14 as=3.0336e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.4338e-06 sim_w=5.76e-06 m_per_maxw=1.04167 numb_sub_cont=3 nfing=1 $X=33380 $Y=200 $D=22
M14 1 2 1 cpoly_n w=6e-06 l=2e-06 c=7.5402e-14 as=3.0336e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.4338e-06 sim_w=5.76e-06 m_per_maxw=1.04167 numb_sub_cont=3 nfing=1 $X=35900 $Y=200 $D=22
M15 1 2 1 cpoly_n w=6e-06 l=2e-06 c=7.5402e-14 as=3.0336e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.4338e-06 sim_w=5.76e-06 m_per_maxw=1.04167 numb_sub_cont=3 nfing=1 $X=38420 $Y=200 $D=22
M16 1 2 1 cpoly_n w=6e-06 l=2e-06 c=7.5402e-14 as=3.0336e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.4338e-06 sim_w=5.76e-06 m_per_maxw=1.04167 numb_sub_cont=3 nfing=1 $X=40940 $Y=200 $D=22
M17 1 2 1 cpoly_n w=6e-06 l=2e-06 c=7.5402e-14 as=3.0336e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.4338e-06 sim_w=5.76e-06 m_per_maxw=1.04167 numb_sub_cont=3 nfing=1 $X=43460 $Y=200 $D=22
M18 1 2 1 cpoly_n w=6e-06 l=2e-06 c=7.5402e-14 as=3.0336e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.4338e-06 sim_w=5.76e-06 m_per_maxw=1.04167 numb_sub_cont=3 nfing=1 $X=45980 $Y=200 $D=22
M19 1 2 1 cpoly_n w=6e-06 l=2e-06 c=7.5402e-14 as=2.4e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.4338e-06 sim_w=5.76e-06 m_per_maxw=1.04167 numb_sub_cont=3 nfing=1 $X=48500 $Y=200 $D=22
.ENDS
***************************************
.SUBCKT Fill_Bit_512x16 gnd! vdd! 7 8 9 10
** N=22 EP=6 IP=52 FDC=214
*.SEEDPROM
M0 12 11 gnd! gnd! nmos_a L=3.8e-07 W=4.8e-07 AD=9.258e-13 AS=2.496e-13 PD=1.06e-06 PS=5.3e-07 w_cont=5.8e-07 nfing=1 source_num=2 $X=12160 $Y=60720 $D=1
M1 14 13 gnd! gnd! nmos_a L=3.8e-07 W=4.8e-07 AD=9.258e-13 AS=1.92e-13 PD=1.06e-06 PS=5.3e-07 w_cont=5.8e-07 nfing=1 source_num=2 $X=24960 $Y=60720 $D=1
M2 16 15 gnd! gnd! nmos_a L=3.8e-07 W=4.8e-07 AD=9.258e-13 AS=2.496e-13 PD=1.06e-06 PS=5.3e-07 w_cont=5.8e-07 nfing=1 source_num=2 $X=13060 $Y=60720 $D=1
M3 18 17 gnd! gnd! nmos_a L=3.8e-07 W=4.8e-07 AD=9.258e-13 AS=2.496e-13 PD=1.06e-06 PS=5.3e-07 w_cont=5.8e-07 nfing=1 source_num=2 $X=38400 $Y=60720 $D=1
M4 20 19 gnd! gnd! nmos_a L=3.8e-07 W=4.8e-07 AD=9.258e-13 AS=1.92e-13 PD=1.06e-06 PS=5.3e-07 w_cont=5.8e-07 nfing=1 source_num=2 $X=26500 $Y=60720 $D=1
M5 22 21 gnd! gnd! nmos_a L=3.8e-07 W=4.8e-07 AD=9.258e-13 AS=2.496e-13 PD=1.06e-06 PS=5.3e-07 w_cont=5.8e-07 nfing=1 source_num=2 $X=39300 $Y=60720 $D=1
X6 gnd! vdd! 11 12 7 8 ICV_29 $T=3200 63000 0 180 $X=-360 $Y=56760
X7 gnd! vdd! 13 14 15 16 ICV_29 $T=16000 63000 0 180 $X=12440 $Y=56760
X8 gnd! vdd! 17 18 19 20 ICV_29 $T=29440 63000 0 180 $X=25880 $Y=56760
X9 gnd! vdd! 9 10 21 22 ICV_29 $T=42240 63000 0 180 $X=38680 $Y=56760
X10 gnd! vdd! cpoly_p_CDNS_58870478665103 $T=460 74440 0 0 $X=460 $Y=74440
X11 gnd! vdd! cpoly_p_CDNS_58870478665103 $T=460 93660 0 0 $X=460 $Y=93660
X12 gnd! vdd! cpoly_p_CDNS_58870478665103 $T=460 112880 0 0 $X=460 $Y=112880
X13 vdd! gnd! cpoly_n_CDNS_58870478665102 $T=51580 65080 1 180 $X=460 $Y=65080
X14 vdd! gnd! cpoly_n_CDNS_58870478665102 $T=51580 84300 1 180 $X=460 $Y=84300
X15 vdd! gnd! cpoly_n_CDNS_58870478665102 $T=51580 103520 1 180 $X=460 $Y=103520
.ENDS
***************************************
.SUBCKT cpoly_p_CDNS_58870478665100 1 2
** N=2 EP=2 IP=0 FDC=10
M0 1 2 1 cpoly_p w=6e-06 l=2e-06 c=8.0712e-14 as=1.68e-13 ad=7.488e-13 ps=1.44e-06 pd=1.13684e-06 sim_w=2.88e-06 m_per_maxw=2.08333 numb_sub_cont=4 nfing=1 $X=620 $Y=200 $D=21
M1 1 2 1 cpoly_p w=6e-06 l=2e-06 c=8.0712e-14 as=2.1408e-13 ad=7.488e-13 ps=1.44e-06 pd=1.13684e-06 sim_w=2.88e-06 m_per_maxw=2.08333 numb_sub_cont=4 nfing=1 $X=3140 $Y=200 $D=21
M2 1 2 1 cpoly_p w=6e-06 l=2e-06 c=8.0712e-14 as=2.1408e-13 ad=7.488e-13 ps=1.44e-06 pd=1.13684e-06 sim_w=2.88e-06 m_per_maxw=2.08333 numb_sub_cont=4 nfing=1 $X=5660 $Y=200 $D=21
M3 1 2 1 cpoly_p w=6e-06 l=2e-06 c=8.0712e-14 as=2.1408e-13 ad=7.488e-13 ps=1.44e-06 pd=1.13684e-06 sim_w=2.88e-06 m_per_maxw=2.08333 numb_sub_cont=4 nfing=1 $X=8180 $Y=200 $D=21
M4 1 2 1 cpoly_p w=6e-06 l=2e-06 c=8.0712e-14 as=2.1408e-13 ad=7.488e-13 ps=1.44e-06 pd=1.13684e-06 sim_w=2.88e-06 m_per_maxw=2.08333 numb_sub_cont=4 nfing=1 $X=10700 $Y=200 $D=21
M5 1 2 1 cpoly_p w=6e-06 l=2e-06 c=8.0712e-14 as=2.1408e-13 ad=7.488e-13 ps=1.44e-06 pd=1.13684e-06 sim_w=2.88e-06 m_per_maxw=2.08333 numb_sub_cont=4 nfing=1 $X=13220 $Y=200 $D=21
M6 1 2 1 cpoly_p w=6e-06 l=2e-06 c=8.0712e-14 as=2.1408e-13 ad=7.488e-13 ps=1.44e-06 pd=1.13684e-06 sim_w=2.88e-06 m_per_maxw=2.08333 numb_sub_cont=4 nfing=1 $X=15740 $Y=200 $D=21
M7 1 2 1 cpoly_p w=6e-06 l=2e-06 c=8.0712e-14 as=2.1408e-13 ad=7.488e-13 ps=1.44e-06 pd=1.13684e-06 sim_w=2.88e-06 m_per_maxw=2.08333 numb_sub_cont=4 nfing=1 $X=18260 $Y=200 $D=21
M8 1 2 1 cpoly_p w=6e-06 l=2e-06 c=8.0712e-14 as=2.1408e-13 ad=7.488e-13 ps=1.44e-06 pd=1.13684e-06 sim_w=2.88e-06 m_per_maxw=2.08333 numb_sub_cont=4 nfing=1 $X=20780 $Y=200 $D=21
M9 1 2 1 cpoly_p w=6e-06 l=2e-06 c=8.0712e-14 as=1.68e-13 ad=7.488e-13 ps=1.44e-06 pd=1.13684e-06 sim_w=2.88e-06 m_per_maxw=2.08333 numb_sub_cont=4 nfing=1 $X=23300 $Y=200 $D=21
.ENDS
***************************************
.SUBCKT cpoly_n_CDNS_58870478665101 1 2
** N=2 EP=2 IP=0 FDC=10
M0 1 2 1 cpoly_n w=6e-06 l=2e-06 c=7.5402e-14 as=2.4e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.4338e-06 sim_w=5.76e-06 m_per_maxw=1.04167 numb_sub_cont=3 nfing=1 $X=620 $Y=200 $D=22
M1 1 2 1 cpoly_n w=6e-06 l=2e-06 c=7.5402e-14 as=3.0336e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.4338e-06 sim_w=5.76e-06 m_per_maxw=1.04167 numb_sub_cont=3 nfing=1 $X=3140 $Y=200 $D=22
M2 1 2 1 cpoly_n w=6e-06 l=2e-06 c=7.5402e-14 as=3.0336e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.4338e-06 sim_w=5.76e-06 m_per_maxw=1.04167 numb_sub_cont=3 nfing=1 $X=5660 $Y=200 $D=22
M3 1 2 1 cpoly_n w=6e-06 l=2e-06 c=7.5402e-14 as=3.0336e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.4338e-06 sim_w=5.76e-06 m_per_maxw=1.04167 numb_sub_cont=3 nfing=1 $X=8180 $Y=200 $D=22
M4 1 2 1 cpoly_n w=6e-06 l=2e-06 c=7.5402e-14 as=3.0336e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.4338e-06 sim_w=5.76e-06 m_per_maxw=1.04167 numb_sub_cont=3 nfing=1 $X=10700 $Y=200 $D=22
M5 1 2 1 cpoly_n w=6e-06 l=2e-06 c=7.5402e-14 as=3.0336e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.4338e-06 sim_w=5.76e-06 m_per_maxw=1.04167 numb_sub_cont=3 nfing=1 $X=13220 $Y=200 $D=22
M6 1 2 1 cpoly_n w=6e-06 l=2e-06 c=7.5402e-14 as=3.0336e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.4338e-06 sim_w=5.76e-06 m_per_maxw=1.04167 numb_sub_cont=3 nfing=1 $X=15740 $Y=200 $D=22
M7 1 2 1 cpoly_n w=6e-06 l=2e-06 c=7.5402e-14 as=3.0336e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.4338e-06 sim_w=5.76e-06 m_per_maxw=1.04167 numb_sub_cont=3 nfing=1 $X=18260 $Y=200 $D=22
M8 1 2 1 cpoly_n w=6e-06 l=2e-06 c=7.5402e-14 as=3.0336e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.4338e-06 sim_w=5.76e-06 m_per_maxw=1.04167 numb_sub_cont=3 nfing=1 $X=20780 $Y=200 $D=22
M9 1 2 1 cpoly_n w=6e-06 l=2e-06 c=7.5402e-14 as=2.4e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.4338e-06 sim_w=5.76e-06 m_per_maxw=1.04167 numb_sub_cont=3 nfing=1 $X=23300 $Y=200 $D=22
.ENDS
***************************************
.SUBCKT Fill_Block_8Kx8 gnd! vdd!
** N=41 EP=2 IP=92 FDC=1788
M0 11 10 gnd! gnd! nmos_a L=3.8e-07 W=4.8e-07 AD=9.258e-13 AS=1.92e-13 PD=1.06e-06 PS=5.3e-07 w_cont=5.8e-07 nfing=1 source_num=2 $X=260 $Y=60820 $D=1
M1 13 12 gnd! gnd! nmos_a L=3.8e-07 W=4.8e-07 AD=9.258e-13 AS=2.496e-13 PD=1.06e-06 PS=5.3e-07 w_cont=5.8e-07 nfing=1 source_num=2 $X=51200 $Y=60820 $D=1
M2 15 14 gnd! gnd! nmos_a L=3.8e-07 W=4.8e-07 AD=9.258e-13 AS=2.496e-13 PD=1.06e-06 PS=5.3e-07 w_cont=5.8e-07 nfing=1 source_num=2 $X=52100 $Y=60820 $D=1
M3 17 16 gnd! gnd! nmos_a L=3.8e-07 W=4.8e-07 AD=9.258e-13 AS=2.496e-13 PD=1.06e-06 PS=5.3e-07 w_cont=5.8e-07 nfing=1 source_num=2 $X=103040 $Y=60820 $D=1
M4 19 18 gnd! gnd! nmos_a L=3.8e-07 W=4.8e-07 AD=9.258e-13 AS=2.496e-13 PD=1.06e-06 PS=5.3e-07 w_cont=5.8e-07 nfing=1 source_num=2 $X=103940 $Y=60820 $D=1
M5 21 20 gnd! gnd! nmos_a L=3.8e-07 W=4.8e-07 AD=9.258e-13 AS=2.496e-13 PD=1.06e-06 PS=5.3e-07 w_cont=5.8e-07 nfing=1 source_num=2 $X=154880 $Y=60820 $D=1
M6 23 22 gnd! gnd! nmos_a L=3.8e-07 W=4.8e-07 AD=9.258e-13 AS=2.496e-13 PD=1.06e-06 PS=5.3e-07 w_cont=5.8e-07 nfing=1 source_num=2 $X=155780 $Y=60820 $D=1
M7 25 24 gnd! gnd! nmos_a L=3.8e-07 W=4.8e-07 AD=9.258e-13 AS=1.92e-13 PD=1.06e-06 PS=5.3e-07 w_cont=5.8e-07 nfing=1 source_num=2 $X=206720 $Y=60820 $D=1
M8 27 26 gnd! gnd! nmos_a L=3.8e-07 W=4.8e-07 AD=9.258e-13 AS=1.92e-13 PD=1.06e-06 PS=5.3e-07 w_cont=5.8e-07 nfing=1 source_num=2 $X=232740 $Y=60820 $D=1
M9 29 28 gnd! gnd! nmos_a L=3.8e-07 W=4.8e-07 AD=9.258e-13 AS=2.496e-13 PD=1.06e-06 PS=5.3e-07 w_cont=5.8e-07 nfing=1 source_num=2 $X=283680 $Y=60820 $D=1
M10 31 30 gnd! gnd! nmos_a L=3.8e-07 W=4.8e-07 AD=9.258e-13 AS=2.496e-13 PD=1.06e-06 PS=5.3e-07 w_cont=5.8e-07 nfing=1 source_num=2 $X=284580 $Y=60820 $D=1
M11 33 32 gnd! gnd! nmos_a L=3.8e-07 W=4.8e-07 AD=9.258e-13 AS=2.496e-13 PD=1.06e-06 PS=5.3e-07 w_cont=5.8e-07 nfing=1 source_num=2 $X=335520 $Y=60820 $D=1
M12 35 34 gnd! gnd! nmos_a L=3.8e-07 W=4.8e-07 AD=9.258e-13 AS=2.496e-13 PD=1.06e-06 PS=5.3e-07 w_cont=5.8e-07 nfing=1 source_num=2 $X=336420 $Y=60820 $D=1
M13 37 36 gnd! gnd! nmos_a L=3.8e-07 W=4.8e-07 AD=9.258e-13 AS=2.496e-13 PD=1.06e-06 PS=5.3e-07 w_cont=5.8e-07 nfing=1 source_num=2 $X=387360 $Y=60820 $D=1
M14 39 38 gnd! gnd! nmos_a L=3.8e-07 W=4.8e-07 AD=9.258e-13 AS=2.496e-13 PD=1.06e-06 PS=5.3e-07 w_cont=5.8e-07 nfing=1 source_num=2 $X=388260 $Y=60820 $D=1
M15 41 40 gnd! gnd! nmos_a L=3.8e-07 W=4.8e-07 AD=9.258e-13 AS=1.92e-13 PD=1.06e-06 PS=5.3e-07 w_cont=5.8e-07 nfing=1 source_num=2 $X=439200 $Y=60820 $D=1
X16 gnd! vdd! 10 11 12 13 Fill_Bit_512x16 $T=0 122600 1 0 $X=-360 $Y=-320
X17 gnd! vdd! 14 15 16 17 Fill_Bit_512x16 $T=51840 122600 1 0 $X=51480 $Y=-320
X18 gnd! vdd! 18 19 20 21 Fill_Bit_512x16 $T=103680 122600 1 0 $X=103320 $Y=-320
X19 gnd! vdd! 22 23 24 25 Fill_Bit_512x16 $T=155520 122600 1 0 $X=155160 $Y=-320
X20 gnd! vdd! 26 27 28 29 Fill_Bit_512x16 $T=232480 122600 1 0 $X=232120 $Y=-320
X21 gnd! vdd! 30 31 32 33 Fill_Bit_512x16 $T=284320 122600 1 0 $X=283960 $Y=-320
X22 gnd! vdd! 34 35 36 37 Fill_Bit_512x16 $T=336160 122600 1 0 $X=335800 $Y=-320
X23 gnd! vdd! 38 39 40 41 Fill_Bit_512x16 $T=388000 122600 1 0 $X=387640 $Y=-320
X24 gnd! vdd! cpoly_p_CDNS_58870478665100 $T=232980 9720 0 180 $X=207060 $Y=1720
X25 gnd! vdd! cpoly_p_CDNS_58870478665100 $T=232980 28940 0 180 $X=207060 $Y=20940
X26 gnd! vdd! cpoly_p_CDNS_58870478665100 $T=232980 48160 0 180 $X=207060 $Y=40160
X27 vdd! gnd! cpoly_n_CDNS_58870478665101 $T=207060 19080 1 0 $X=207060 $Y=11580
X28 vdd! gnd! cpoly_n_CDNS_58870478665101 $T=207060 38300 1 0 $X=207060 $Y=30800
X29 vdd! gnd! cpoly_n_CDNS_58870478665101 $T=207060 57520 1 0 $X=207060 $Y=50020
.ENDS
***************************************
.SUBCKT nmos_a_CDNS_5887047866586 1 2 3
** N=3 EP=3 IP=0 FDC=3
M0 2 3 1 1 nmos_a L=2.4e-07 W=3.6e-06 AD=1.0816e-12 AS=1.44e-12 PD=2.08e-06 PS=2.08e-06 w_cont=1.6e-06 nfing=1 source_num=2 $X=620 $Y=200 $D=1
M1 2 3 1 1 nmos_a L=2.4e-07 W=3.6e-06 AD=1.0816e-12 AS=9.36e-13 PD=2.08e-06 PS=2.08e-06 w_cont=1.6e-06 nfing=1 source_num=2 $X=1380 $Y=200 $D=1
M2 2 3 1 1 nmos_a L=2.4e-07 W=3.6e-06 AD=1.664e-12 AS=9.36e-13 PD=4.16e-06 PS=2.08e-06 w_cont=1.6e-06 nfing=1 source_num=2 $X=2140 $Y=200 $D=1
.ENDS
***************************************
.SUBCKT pmos_a_CDNS_5887047866522
** N=3 EP=0 IP=0 FDC=0
*.SEEDPROM
.ENDS
***************************************
.SUBCKT pmos_a_CDNS_5887047866592 1 2 3 4
** N=4 EP=4 IP=0 FDC=4
M0 2 3 1 1 pmos_a L=2.4e-07 W=4e-06 AD=1.196e-12 AS=1.4e-13 PD=2.3e-06 PS=2.3e-06 w_cont=6e-07 nfing=1 mmm=1 $X=620 $Y=200 $D=5
M1 2 3 1 1 pmos_a L=2.4e-07 W=4e-06 AD=1.196e-12 AS=1.76e-13 PD=2.3e-06 PS=2.3e-06 w_cont=6e-07 nfing=1 mmm=1 $X=1380 $Y=200 $D=5
M2 2 4 1 1 pmos_a L=2.4e-07 W=4e-06 AD=1.196e-12 AS=1.76e-13 PD=2.3e-06 PS=2.3e-06 w_cont=6e-07 nfing=1 mmm=1 $X=2140 $Y=200 $D=5
M3 2 4 1 1 pmos_a L=2.4e-07 W=4e-06 AD=1.196e-12 AS=1.4e-13 PD=2.3e-06 PS=2.3e-06 w_cont=6e-07 nfing=1 mmm=1 $X=2900 $Y=200 $D=5
.ENDS
***************************************
.SUBCKT nmos_io_a_CDNS_5887047866594 1 2 3
** N=3 EP=3 IP=0 FDC=1
M0 2 3 1 1 nmos_io_a L=2.8e-07 W=4.8e-06 AD=7.5348e-12 AS=2.664e-13 PD=4.14e-06 PS=2.07e-06 w_cont=2.1e-06 nfing=1 $X=620 $Y=200 $D=0
.ENDS
***************************************
.SUBCKT dn_CDNS_5887047866588 1 2
** N=2 EP=2 IP=0 FDC=1
D0 2 1 dn PJ=4e-06 m=1 $X=-460 $Y=0 $D=9
.ENDS
***************************************
.SUBCKT pmos_io_a_CDNS_5887047866595 1 2 3
** N=3 EP=3 IP=0 FDC=1
M0 2 3 1 1 pmos_io_a L=2.8e-07 W=9e-06 AD=1.17645e-11 AS=1.696e-13 PD=6.464e-06 PS=3.232e-06 w_cont=1.1e-06 nfing=1 $X=620 $Y=200 $D=4
.ENDS
***************************************
.SUBCKT cpoly_n_CDNS_5887047866515 1 2
** N=2 EP=2 IP=0 FDC=6
M0 1 2 1 cpoly_n w=6e-06 l=2e-06 c=7.5402e-14 as=2.4e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.4338e-06 sim_w=5.76e-06 m_per_maxw=1.04167 numb_sub_cont=3 nfing=1 $X=620 $Y=200 $D=22
M1 1 2 1 cpoly_n w=6e-06 l=2e-06 c=7.5402e-14 as=3.0336e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.4338e-06 sim_w=5.76e-06 m_per_maxw=1.04167 numb_sub_cont=3 nfing=1 $X=3140 $Y=200 $D=22
M2 1 2 1 cpoly_n w=6e-06 l=2e-06 c=7.5402e-14 as=3.0336e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.4338e-06 sim_w=5.76e-06 m_per_maxw=1.04167 numb_sub_cont=3 nfing=1 $X=5660 $Y=200 $D=22
M3 1 2 1 cpoly_n w=6e-06 l=2e-06 c=7.5402e-14 as=3.0336e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.4338e-06 sim_w=5.76e-06 m_per_maxw=1.04167 numb_sub_cont=3 nfing=1 $X=8180 $Y=200 $D=22
M4 1 2 1 cpoly_n w=6e-06 l=2e-06 c=7.5402e-14 as=3.0336e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.4338e-06 sim_w=5.76e-06 m_per_maxw=1.04167 numb_sub_cont=3 nfing=1 $X=10700 $Y=200 $D=22
M5 1 2 1 cpoly_n w=6e-06 l=2e-06 c=7.5402e-14 as=2.4e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.4338e-06 sim_w=5.76e-06 m_per_maxw=1.04167 numb_sub_cont=3 nfing=1 $X=13220 $Y=200 $D=22
.ENDS
***************************************
.SUBCKT nmos_a_CDNS_5887047866587
** N=3 EP=0 IP=0 FDC=0
*.SEEDPROM
.ENDS
***************************************
.SUBCKT PADIO nWE GND_PAD VDD_PAD gnd! vdd! DIO DI DO nOE
** N=36 EP=9 IP=412 FDC=293
M0 15 36 gnd! gnd! nmos_a L=2.4e-07 W=4.8e-07 AD=4.32e-13 AS=2.496e-13 PD=1.08e-06 PS=5.4e-07 w_cont=6e-07 nfing=1 source_num=2 $X=10440 $Y=326780 $D=1
M1 19 21 gnd! gnd! nmos_a L=2.4e-07 W=4.8e-07 AD=4.32e-13 AS=2.496e-13 PD=1.08e-06 PS=5.4e-07 w_cont=6e-07 nfing=1 source_num=2 $X=11200 $Y=326780 $D=1
M2 13 28 26 26 nmos_a L=2.4e-07 W=2.4e-06 AD=1.4e-12 AS=9.6e-13 PD=3.5e-06 PS=1.75e-06 w_cont=1.1e-06 nfing=1 source_num=2 $X=76440 $Y=317040 $D=1
M3 33 34 35 35 nmos_a L=2.4e-07 W=2.4e-06 AD=1.4e-12 AS=9.6e-13 PD=3.5e-06 PS=1.75e-06 w_cont=1.1e-06 nfing=1 source_num=2 $X=91660 $Y=332540 $D=1
M4 35 31 gnd! gnd! nmos_a L=2.4e-07 W=2.4e-06 AD=1.4e-12 AS=9.6e-13 PD=3.5e-06 PS=1.75e-06 w_cont=1.1e-06 nfing=1 source_num=2 $X=93100 $Y=332540 $D=1
M5 30 31 gnd! gnd! nmos_a L=2.4e-07 W=1.2e-06 AD=7.2e-13 AS=4.8e-13 PD=1.8e-06 PS=9e-07 w_cont=6e-07 nfing=1 source_num=2 $X=83340 $Y=330860 $D=1
M6 34 DO gnd! gnd! nmos_a L=2.4e-07 W=1.2e-06 AD=7.2e-13 AS=4.8e-13 PD=1.8e-06 PS=9e-07 w_cont=6e-07 nfing=1 source_num=2 $X=83440 $Y=335820 $D=1
M7 34 DO gnd! gnd! nmos_a L=2.4e-07 W=1.2e-06 AD=7.2e-13 AS=4.8e-13 PD=1.8e-06 PS=9e-07 w_cont=6e-07 nfing=1 source_num=2 $X=84880 $Y=335820 $D=1
M8 31 nOE gnd! gnd! nmos_a L=2.4e-07 W=1.2e-06 AD=7.2e-13 AS=4.8e-13 PD=1.8e-06 PS=9e-07 w_cont=6e-07 nfing=1 source_num=2 $X=85580 $Y=330520 $D=1
M9 DI 17 gnd! gnd! nmos_a L=2.4e-07 W=4.8e-07 AD=4.32e-13 AS=1.92e-13 PD=1.08e-06 PS=5.4e-07 w_cont=6e-07 nfing=1 source_num=2 $X=8960 $Y=328820 $D=1
M10 17 22 15 15 nmos_a L=2.4e-07 W=4.8e-07 AD=2.808e-13 AS=1.92e-13 PD=5.4e-07 PS=5.4e-07 w_cont=6e-07 nfing=1 source_num=2 $X=10440 $Y=328820 $D=1
M11 17 20 19 19 nmos_a L=2.4e-07 W=4.8e-07 AD=2.808e-13 AS=1.92e-13 PD=5.4e-07 PS=5.4e-07 w_cont=6e-07 nfing=1 source_num=2 $X=11200 $Y=328820 $D=1
M12 21 24 gnd! gnd! nmos_a L=2.4e-07 W=4.8e-07 AD=4.32e-13 AS=1.92e-13 PD=1.08e-06 PS=5.4e-07 w_cont=6e-07 nfing=1 source_num=2 $X=13180 $Y=337900 $D=1
M13 20 22 gnd! gnd! nmos_a L=2.4e-07 W=4.8e-07 AD=4.32e-13 AS=1.92e-13 PD=1.08e-06 PS=5.4e-07 w_cont=6e-07 nfing=1 source_num=2 $X=13680 $Y=329220 $D=1
M14 25 21 gnd! gnd! nmos_a L=2.4e-07 W=4.8e-07 AD=4.32e-13 AS=2.496e-13 PD=1.08e-06 PS=5.4e-07 w_cont=6e-07 nfing=1 source_num=2 $X=14520 $Y=340560 $D=1
M15 22 nWE gnd! gnd! nmos_a L=2.4e-07 W=4.8e-07 AD=4.32e-13 AS=1.92e-13 PD=1.08e-06 PS=5.4e-07 w_cont=6e-07 nfing=1 source_num=2 $X=15120 $Y=329220 $D=1
M16 24 DI 25 25 nmos_a L=4.8e-07 W=4.8e-07 AD=4.32e-13 AS=1.92e-13 PD=1.08e-06 PS=5.4e-07 w_cont=6e-07 nfing=1 source_num=2 $X=15280 $Y=338600 $D=1
M17 25 DI gnd! gnd! nmos_a L=4.8e-07 W=4.8e-07 AD=4.32e-13 AS=2.496e-13 PD=1.08e-06 PS=5.4e-07 w_cont=6e-07 nfing=1 source_num=2 $X=15280 $Y=340560 $D=1
M18 16 21 vdd! vdd! pmos_a L=2.4e-07 W=4.8e-07 AD=4.32e-13 AS=1.584e-13 PD=1.08e-06 PS=5.4e-07 w_cont=6e-07 nfing=1 mmm=1 $X=10440 $Y=334320 $D=5
M19 18 36 vdd! vdd! pmos_a L=2.4e-07 W=4.8e-07 AD=4.32e-13 AS=1.584e-13 PD=1.08e-06 PS=5.4e-07 w_cont=6e-07 nfing=1 mmm=1 $X=11200 $Y=334320 $D=5
M20 13 28 vdd! vdd! pmos_a L=2.4e-07 W=4e-06 AD=1.84e-12 AS=1.76e-13 PD=4.6e-06 PS=2.3e-06 w_cont=6e-07 nfing=1 mmm=1 $X=71960 $Y=317040 $D=5
M21 13 28 vdd! vdd! pmos_a L=2.4e-07 W=4e-06 AD=1.196e-12 AS=1.76e-13 PD=2.3e-06 PS=2.3e-06 w_cont=6e-07 nfing=1 mmm=1 $X=72720 $Y=317040 $D=5
M22 13 28 vdd! vdd! pmos_a L=2.4e-07 W=4e-06 AD=1.196e-12 AS=1.76e-13 PD=2.3e-06 PS=2.3e-06 w_cont=6e-07 nfing=1 mmm=1 $X=73480 $Y=317040 $D=5
M23 13 28 vdd! vdd! pmos_a L=2.4e-07 W=4e-06 AD=1.196e-12 AS=1.76e-13 PD=2.3e-06 PS=2.3e-06 w_cont=6e-07 nfing=1 mmm=1 $X=74240 $Y=317040 $D=5
M24 13 28 vdd! vdd! pmos_a L=2.4e-07 W=4e-06 AD=1.196e-12 AS=1.4e-13 PD=2.3e-06 PS=2.3e-06 w_cont=6e-07 nfing=1 mmm=1 $X=75000 $Y=317040 $D=5
M25 30 31 vdd! vdd! pmos_a L=2.4e-07 W=2e-06 AD=1.04e-12 AS=1.3e-13 PD=2.6e-06 PS=1.3e-06 w_cont=6e-07 nfing=1 mmm=1 $X=83300 $Y=326420 $D=5
M26 34 DO vdd! vdd! pmos_a L=2.4e-07 W=2e-06 AD=1.04e-12 AS=1.3e-13 PD=2.6e-06 PS=1.3e-06 w_cont=6e-07 nfing=1 mmm=1 $X=83440 $Y=338560 $D=5
M27 34 DO vdd! vdd! pmos_a L=2.4e-07 W=2e-06 AD=1.04e-12 AS=1.3e-13 PD=2.6e-06 PS=1.3e-06 w_cont=6e-07 nfing=1 mmm=1 $X=84880 $Y=338560 $D=5
M28 31 nOE vdd! vdd! pmos_a L=2.4e-07 W=2e-06 AD=1.04e-12 AS=1.3e-13 PD=2.6e-06 PS=1.3e-06 w_cont=6e-07 nfing=1 mmm=1 $X=85580 $Y=326420 $D=5
M29 DI 17 vdd! vdd! pmos_a L=2.4e-07 W=1e-06 AD=6.4e-13 AS=1.25e-13 PD=1.6e-06 PS=8e-07 w_cont=6e-07 nfing=1 mmm=1 $X=9000 $Y=331460 $D=5
M30 21 24 vdd! vdd! pmos_a L=2.4e-07 W=1e-06 AD=6.4e-13 AS=1.61e-13 PD=1.6e-06 PS=8e-07 w_cont=6e-07 nfing=1 mmm=1 $X=13320 $Y=334760 $D=5
M31 20 22 vdd! vdd! pmos_a L=2.4e-07 W=1e-06 AD=6.4e-13 AS=1.25e-13 PD=1.6e-06 PS=8e-07 w_cont=6e-07 nfing=1 mmm=1 $X=13680 $Y=331560 $D=5
M32 23 21 vdd! vdd! pmos_a L=2.4e-07 W=1e-06 AD=6.4e-13 AS=1.61e-13 PD=1.6e-06 PS=8e-07 w_cont=6e-07 nfing=1 mmm=1 $X=14080 $Y=334760 $D=5
M33 22 nWE vdd! vdd! pmos_a L=2.4e-07 W=1e-06 AD=6.4e-13 AS=1.25e-13 PD=1.6e-06 PS=8e-07 w_cont=6e-07 nfing=1 mmm=1 $X=15120 $Y=332060 $D=5
M34 17 22 16 16 pmos_a L=2.4e-07 W=4.8e-07 AD=2.808e-13 AS=1.224e-13 PD=5.4e-07 PS=5.4e-07 w_cont=6e-07 nfing=1 mmm=1 $X=10440 $Y=331980 $D=5
M35 17 20 18 18 pmos_a L=2.4e-07 W=4.8e-07 AD=2.808e-13 AS=1.224e-13 PD=5.4e-07 PS=5.4e-07 w_cont=6e-07 nfing=1 mmm=1 $X=11200 $Y=331980 $D=5
M36 23 DI vdd! vdd! pmos_a L=2.4e-07 W=4.8e-07 AD=4.32e-13 AS=1.224e-13 PD=1.08e-06 PS=5.4e-07 w_cont=6e-07 nfing=1 mmm=1 $X=15520 $Y=334760 $D=5
M37 24 DI 23 23 pmos_a L=2.4e-07 W=4.8e-07 AD=4.32e-13 AS=1.224e-13 PD=1.08e-06 PS=5.4e-07 w_cont=6e-07 nfing=1 mmm=1 $X=15520 $Y=336620 $D=5
M38 32 29 vdd! vdd! pmos_a L=2.4e-07 W=4e-06 AD=1.84e-12 AS=1.4e-13 PD=4.6e-06 PS=2.3e-06 w_cont=6e-07 nfing=1 mmm=1 $X=88860 $Y=317040 $D=5
M39 14 33 32 32 pmos_a L=2.4e-07 W=4e-06 AD=1.84e-12 AS=1.4e-13 PD=4.6e-06 PS=2.3e-06 w_cont=6e-07 nfing=1 mmm=1 $X=90300 $Y=317040 $D=5
M40 gnd! 24 gnd! cpoly_p w=6e-06 l=2e-06 c=8.0712e-14 as=2.1408e-13 ad=1.152e-12 ps=1.44e-06 pd=2.27368e-06 sim_w=2.88e-06 m_per_maxw=2.08333 numb_sub_cont=4 nfing=1 $X=8180 $Y=317980 $D=21
M41 gnd! 24 gnd! cpoly_p w=6e-06 l=2e-06 c=8.0712e-14 as=2.1408e-13 ad=7.488e-13 ps=1.44e-06 pd=1.13684e-06 sim_w=2.88e-06 m_per_maxw=2.08333 numb_sub_cont=4 nfing=1 $X=10700 $Y=317980 $D=21
M42 gnd! 24 gnd! cpoly_p w=6e-06 l=2e-06 c=8.0712e-14 as=1.68e-13 ad=7.488e-13 ps=1.44e-06 pd=1.13684e-06 sim_w=2.88e-06 m_per_maxw=2.08333 numb_sub_cont=4 nfing=1 $X=13220 $Y=317980 $D=21
M43 gnd! vdd! gnd! cpoly_p w=6e-06 l=2e-06 c=8.0712e-14 as=1.68e-13 ad=7.488e-13 ps=1.44e-06 pd=1.13684e-06 sim_w=2.88e-06 m_per_maxw=2.08333 numb_sub_cont=4 nfing=1 $X=17000 $Y=317980 $D=21
M44 gnd! vdd! gnd! cpoly_p w=6e-06 l=2e-06 c=8.0712e-14 as=2.1408e-13 ad=7.488e-13 ps=1.44e-06 pd=1.13684e-06 sim_w=2.88e-06 m_per_maxw=2.08333 numb_sub_cont=4 nfing=1 $X=19520 $Y=317980 $D=21
M45 gnd! vdd! gnd! cpoly_p w=6e-06 l=2e-06 c=8.0712e-14 as=2.1408e-13 ad=7.488e-13 ps=1.44e-06 pd=1.13684e-06 sim_w=2.88e-06 m_per_maxw=2.08333 numb_sub_cont=4 nfing=1 $X=22040 $Y=317980 $D=21
M46 gnd! vdd! gnd! cpoly_p w=6e-06 l=2e-06 c=8.0712e-14 as=2.1408e-13 ad=7.488e-13 ps=1.44e-06 pd=1.13684e-06 sim_w=2.88e-06 m_per_maxw=2.08333 numb_sub_cont=4 nfing=1 $X=24560 $Y=317980 $D=21
M47 gnd! vdd! gnd! cpoly_p w=6e-06 l=2e-06 c=8.0712e-14 as=2.1408e-13 ad=7.488e-13 ps=1.44e-06 pd=1.13684e-06 sim_w=2.88e-06 m_per_maxw=2.08333 numb_sub_cont=4 nfing=1 $X=27080 $Y=317980 $D=21
M48 gnd! vdd! gnd! cpoly_p w=6e-06 l=2e-06 c=8.0712e-14 as=2.1408e-13 ad=7.488e-13 ps=1.44e-06 pd=1.13684e-06 sim_w=2.88e-06 m_per_maxw=2.08333 numb_sub_cont=4 nfing=1 $X=29600 $Y=317980 $D=21
M49 gnd! vdd! gnd! cpoly_p w=6e-06 l=2e-06 c=8.0712e-14 as=2.1408e-13 ad=7.488e-13 ps=1.44e-06 pd=1.13684e-06 sim_w=2.88e-06 m_per_maxw=2.08333 numb_sub_cont=4 nfing=1 $X=32120 $Y=317980 $D=21
M50 gnd! vdd! gnd! cpoly_p w=6e-06 l=2e-06 c=8.0712e-14 as=2.1408e-13 ad=7.488e-13 ps=1.44e-06 pd=1.13684e-06 sim_w=2.88e-06 m_per_maxw=2.08333 numb_sub_cont=4 nfing=1 $X=34640 $Y=317980 $D=21
M51 gnd! vdd! gnd! cpoly_p w=6e-06 l=2e-06 c=8.0712e-14 as=2.1408e-13 ad=7.488e-13 ps=1.44e-06 pd=1.13684e-06 sim_w=2.88e-06 m_per_maxw=2.08333 numb_sub_cont=4 nfing=1 $X=37160 $Y=317980 $D=21
M52 gnd! vdd! gnd! cpoly_p w=6e-06 l=2e-06 c=8.0712e-14 as=2.1408e-13 ad=7.488e-13 ps=1.44e-06 pd=1.13684e-06 sim_w=2.88e-06 m_per_maxw=2.08333 numb_sub_cont=4 nfing=1 $X=39680 $Y=317980 $D=21
M53 gnd! vdd! gnd! cpoly_p w=6e-06 l=2e-06 c=8.0712e-14 as=2.1408e-13 ad=7.488e-13 ps=1.44e-06 pd=1.13684e-06 sim_w=2.88e-06 m_per_maxw=2.08333 numb_sub_cont=4 nfing=1 $X=42200 $Y=317980 $D=21
M54 gnd! vdd! gnd! cpoly_p w=6e-06 l=2e-06 c=8.0712e-14 as=2.1408e-13 ad=7.488e-13 ps=1.44e-06 pd=1.13684e-06 sim_w=2.88e-06 m_per_maxw=2.08333 numb_sub_cont=4 nfing=1 $X=44720 $Y=317980 $D=21
M55 gnd! vdd! gnd! cpoly_p w=6e-06 l=2e-06 c=8.0712e-14 as=2.1408e-13 ad=7.488e-13 ps=1.44e-06 pd=1.13684e-06 sim_w=2.88e-06 m_per_maxw=2.08333 numb_sub_cont=4 nfing=1 $X=47240 $Y=317980 $D=21
M56 gnd! vdd! gnd! cpoly_p w=6e-06 l=2e-06 c=8.0712e-14 as=2.1408e-13 ad=7.488e-13 ps=1.44e-06 pd=1.13684e-06 sim_w=2.88e-06 m_per_maxw=2.08333 numb_sub_cont=4 nfing=1 $X=49760 $Y=317980 $D=21
M57 gnd! vdd! gnd! cpoly_p w=6e-06 l=2e-06 c=8.0712e-14 as=2.1408e-13 ad=7.488e-13 ps=1.44e-06 pd=1.13684e-06 sim_w=2.88e-06 m_per_maxw=2.08333 numb_sub_cont=4 nfing=1 $X=52280 $Y=317980 $D=21
M58 gnd! vdd! gnd! cpoly_p w=6e-06 l=2e-06 c=8.0712e-14 as=2.1408e-13 ad=7.488e-13 ps=1.44e-06 pd=1.13684e-06 sim_w=2.88e-06 m_per_maxw=2.08333 numb_sub_cont=4 nfing=1 $X=54800 $Y=317980 $D=21
M59 gnd! vdd! gnd! cpoly_p w=6e-06 l=2e-06 c=8.0712e-14 as=2.1408e-13 ad=7.488e-13 ps=1.44e-06 pd=1.13684e-06 sim_w=2.88e-06 m_per_maxw=2.08333 numb_sub_cont=4 nfing=1 $X=57320 $Y=317980 $D=21
M60 gnd! vdd! gnd! cpoly_p w=6e-06 l=2e-06 c=8.0712e-14 as=2.1408e-13 ad=7.488e-13 ps=1.44e-06 pd=1.13684e-06 sim_w=2.88e-06 m_per_maxw=2.08333 numb_sub_cont=4 nfing=1 $X=59840 $Y=317980 $D=21
M61 gnd! vdd! gnd! cpoly_p w=6e-06 l=2e-06 c=8.0712e-14 as=2.1408e-13 ad=7.488e-13 ps=1.44e-06 pd=1.13684e-06 sim_w=2.88e-06 m_per_maxw=2.08333 numb_sub_cont=4 nfing=1 $X=62360 $Y=317980 $D=21
M62 gnd! vdd! gnd! cpoly_p w=6e-06 l=2e-06 c=8.0712e-14 as=2.1408e-13 ad=7.488e-13 ps=1.44e-06 pd=1.13684e-06 sim_w=2.88e-06 m_per_maxw=2.08333 numb_sub_cont=4 nfing=1 $X=64880 $Y=317980 $D=21
M63 gnd! vdd! gnd! cpoly_p w=6e-06 l=2e-06 c=8.0712e-14 as=2.1408e-13 ad=1.152e-12 ps=1.44e-06 pd=2.27368e-06 sim_w=2.88e-06 m_per_maxw=2.08333 numb_sub_cont=4 nfing=1 $X=67400 $Y=317980 $D=21
M64 gnd! vdd! gnd! cpoly_p w=8.62e-06 l=2e-06 c=1.08536e-13 as=1.21314e-13 ad=1.152e-12 ps=1.44e-06 pd=2.42912e-06 sim_w=2.88e-06 m_per_maxw=2.99306 numb_sub_cont=4 nfing=1 $X=96500 $Y=320700 $D=21
M65 vdd! gnd! vdd! cpoly_n w=6e-06 l=2e-06 c=7.5402e-14 as=2.4e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.4338e-06 sim_w=5.76e-06 m_per_maxw=1.04167 numb_sub_cont=3 nfing=1 $X=1820 $Y=336700 $D=22
M66 vdd! gnd! vdd! cpoly_n w=6e-06 l=2e-06 c=7.5402e-14 as=3.0336e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.4338e-06 sim_w=5.76e-06 m_per_maxw=1.04167 numb_sub_cont=3 nfing=1 $X=4340 $Y=336700 $D=22
M67 vdd! gnd! vdd! cpoly_n w=6e-06 l=2e-06 c=7.5402e-14 as=3.0336e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.4338e-06 sim_w=5.76e-06 m_per_maxw=1.04167 numb_sub_cont=3 nfing=1 $X=6860 $Y=336700 $D=22
M68 vdd! gnd! vdd! cpoly_n w=6e-06 l=2e-06 c=7.5402e-14 as=2.4e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.4338e-06 sim_w=5.76e-06 m_per_maxw=1.04167 numb_sub_cont=3 nfing=1 $X=9380 $Y=336700 $D=22
M69 vdd! gnd! vdd! cpoly_n w=6e-06 l=2e-06 c=7.5402e-14 as=2.4e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.4338e-06 sim_w=5.76e-06 m_per_maxw=1.04167 numb_sub_cont=3 nfing=1 $X=59860 $Y=336700 $D=22
M70 vdd! gnd! vdd! cpoly_n w=6e-06 l=2e-06 c=7.5402e-14 as=3.0336e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.4338e-06 sim_w=5.76e-06 m_per_maxw=1.04167 numb_sub_cont=3 nfing=1 $X=62380 $Y=336700 $D=22
M71 vdd! gnd! vdd! cpoly_n w=6e-06 l=2e-06 c=7.5402e-14 as=3.0336e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.4338e-06 sim_w=5.76e-06 m_per_maxw=1.04167 numb_sub_cont=3 nfing=1 $X=64900 $Y=336700 $D=22
M72 vdd! gnd! vdd! cpoly_n w=6e-06 l=2e-06 c=7.5402e-14 as=3.0336e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.4338e-06 sim_w=5.76e-06 m_per_maxw=1.04167 numb_sub_cont=3 nfing=1 $X=67420 $Y=336700 $D=22
M73 vdd! gnd! vdd! cpoly_n w=6e-06 l=2e-06 c=7.5402e-14 as=3.0336e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.4338e-06 sim_w=5.76e-06 m_per_maxw=1.04167 numb_sub_cont=3 nfing=1 $X=69940 $Y=336700 $D=22
M74 vdd! gnd! vdd! cpoly_n w=6e-06 l=2e-06 c=7.5402e-14 as=3.0336e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.4338e-06 sim_w=5.76e-06 m_per_maxw=1.04167 numb_sub_cont=3 nfing=1 $X=72460 $Y=336700 $D=22
M75 vdd! gnd! vdd! cpoly_n w=6e-06 l=2e-06 c=7.5402e-14 as=3.0336e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.4338e-06 sim_w=5.76e-06 m_per_maxw=1.04167 numb_sub_cont=3 nfing=1 $X=74980 $Y=336700 $D=22
M76 vdd! gnd! vdd! cpoly_n w=6e-06 l=2e-06 c=7.5402e-14 as=3.0336e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.4338e-06 sim_w=5.76e-06 m_per_maxw=1.04167 numb_sub_cont=3 nfing=1 $X=77500 $Y=336700 $D=22
M77 vdd! gnd! vdd! cpoly_n w=6e-06 l=2e-06 c=7.5402e-14 as=3.0336e-13 ad=2.304e-12 ps=2.88e-06 pd=4.86761e-06 sim_w=5.76e-06 m_per_maxw=1.04167 numb_sub_cont=3 nfing=1 $X=80020 $Y=336700 $D=22
M78 vdd! gnd! vdd! cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=1.67141e-13 ad=2.304e-12 ps=2.88e-06 pd=5.14246e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=96280 $Y=333540 $D=22
R79 29 DIO 291.123 L=5e-06 W=2e-06 m=1 $[rnpoly] $X=80300 $Y=315800 $D=18
D80 DIO VDD_PAD dn PJ=0.0002 m=1 $X=4020 $Y=-95300 $D=8
D81 DIO VDD_PAD dn PJ=0.0002 m=1 $X=4020 $Y=114700 $D=8
D82 GND_PAD DIO dn PJ=0.0002 m=1 $X=6340 $Y=-99700 $D=8
D83 GND_PAD DIO dn PJ=0.0002 m=1 $X=6340 $Y=110300 $D=8
D84 DIO VDD_PAD dn PJ=0.0002 m=1 $X=8660 $Y=-95300 $D=8
D85 DIO VDD_PAD dn PJ=0.0002 m=1 $X=8660 $Y=114700 $D=8
D86 GND_PAD DIO dn PJ=0.0001 m=1 $X=10980 $Y=-99700 $D=8
D87 GND_PAD DIO dn PJ=0.0001 m=1 $X=10980 $Y=110300 $D=8
D88 DIO VDD_PAD dn PJ=0.0001 m=1 $X=14160 $Y=4700 $D=8
D89 DIO VDD_PAD dn PJ=0.0001 m=1 $X=14160 $Y=214700 $D=8
D90 GND_PAD DIO dn PJ=0.0002 m=1 $X=16480 $Y=-99700 $D=8
D91 GND_PAD DIO dn PJ=0.0002 m=1 $X=16480 $Y=110300 $D=8
D92 DIO VDD_PAD dn PJ=0.0002 m=1 $X=18800 $Y=-95300 $D=8
D93 DIO VDD_PAD dn PJ=0.0002 m=1 $X=18800 $Y=114700 $D=8
D94 GND_PAD DIO dn PJ=0.0002 m=1 $X=21120 $Y=-99700 $D=8
D95 GND_PAD DIO dn PJ=0.0002 m=1 $X=21120 $Y=110300 $D=8
D96 DIO VDD_PAD dn PJ=0.0002 m=1 $X=23440 $Y=-95300 $D=8
D97 DIO VDD_PAD dn PJ=0.0002 m=1 $X=23440 $Y=114700 $D=8
D98 GND_PAD DIO dn PJ=0.0001 m=1 $X=25760 $Y=-99700 $D=8
D99 GND_PAD DIO dn PJ=0.0001 m=1 $X=25760 $Y=110300 $D=8
D100 DIO VDD_PAD dn PJ=0.0001 m=1 $X=28940 $Y=4700 $D=8
D101 DIO VDD_PAD dn PJ=0.0001 m=1 $X=28940 $Y=214700 $D=8
D102 GND_PAD DIO dn PJ=0.0002 m=1 $X=31260 $Y=-99700 $D=8
D103 GND_PAD DIO dn PJ=0.0002 m=1 $X=31260 $Y=110300 $D=8
D104 DIO VDD_PAD dn PJ=0.0002 m=1 $X=33580 $Y=-95300 $D=8
D105 DIO VDD_PAD dn PJ=0.0002 m=1 $X=33580 $Y=114700 $D=8
D106 GND_PAD DIO dn PJ=0.0002 m=1 $X=35900 $Y=-99700 $D=8
D107 GND_PAD DIO dn PJ=0.0002 m=1 $X=35900 $Y=110300 $D=8
D108 DIO VDD_PAD dn PJ=0.0002 m=1 $X=38220 $Y=-95300 $D=8
D109 DIO VDD_PAD dn PJ=0.0002 m=1 $X=38220 $Y=114700 $D=8
D110 GND_PAD DIO dn PJ=0.0001 m=1 $X=40540 $Y=-99700 $D=8
D111 GND_PAD DIO dn PJ=0.0001 m=1 $X=40540 $Y=110300 $D=8
D112 DIO VDD_PAD dn PJ=0.0001 m=1 $X=43720 $Y=4700 $D=8
D113 DIO VDD_PAD dn PJ=0.0001 m=1 $X=43720 $Y=214700 $D=8
D114 GND_PAD DIO dn PJ=0.0002 m=1 $X=46040 $Y=-99700 $D=8
D115 GND_PAD DIO dn PJ=0.0002 m=1 $X=46040 $Y=110300 $D=8
D116 DIO VDD_PAD dn PJ=0.0002 m=1 $X=48360 $Y=-95300 $D=8
D117 DIO VDD_PAD dn PJ=0.0002 m=1 $X=48360 $Y=114700 $D=8
D118 GND_PAD DIO dn PJ=0.0002 m=1 $X=50680 $Y=-99700 $D=8
D119 GND_PAD DIO dn PJ=0.0002 m=1 $X=50680 $Y=110300 $D=8
D120 DIO VDD_PAD dn PJ=0.0002 m=1 $X=53000 $Y=-95300 $D=8
D121 DIO VDD_PAD dn PJ=0.0002 m=1 $X=53000 $Y=114700 $D=8
D122 GND_PAD DIO dn PJ=0.0001 m=1 $X=55320 $Y=-99700 $D=8
D123 GND_PAD DIO dn PJ=0.0001 m=1 $X=55320 $Y=110300 $D=8
D124 DIO VDD_PAD dn PJ=0.0001 m=1 $X=58500 $Y=4700 $D=8
D125 DIO VDD_PAD dn PJ=0.0001 m=1 $X=58500 $Y=214700 $D=8
D126 GND_PAD DIO dn PJ=0.0002 m=1 $X=60820 $Y=-99700 $D=8
D127 GND_PAD DIO dn PJ=0.0002 m=1 $X=60820 $Y=110300 $D=8
D128 DIO VDD_PAD dn PJ=0.0002 m=1 $X=63140 $Y=-95300 $D=8
D129 DIO VDD_PAD dn PJ=0.0002 m=1 $X=63140 $Y=114700 $D=8
D130 GND_PAD DIO dn PJ=0.0002 m=1 $X=65460 $Y=-99700 $D=8
D131 GND_PAD DIO dn PJ=0.0002 m=1 $X=65460 $Y=110300 $D=8
D132 DIO VDD_PAD dn PJ=0.0002 m=1 $X=67780 $Y=-95300 $D=8
D133 DIO VDD_PAD dn PJ=0.0002 m=1 $X=67780 $Y=114700 $D=8
D134 GND_PAD DIO dn PJ=0.0001 m=1 $X=70100 $Y=-99700 $D=8
D135 GND_PAD DIO dn PJ=0.0001 m=1 $X=70100 $Y=110300 $D=8
D136 DIO VDD_PAD dn PJ=0.0001 m=1 $X=73280 $Y=4700 $D=8
D137 DIO VDD_PAD dn PJ=0.0001 m=1 $X=73280 $Y=214700 $D=8
D138 GND_PAD DIO dn PJ=0.0002 m=1 $X=75600 $Y=-99700 $D=8
D139 GND_PAD DIO dn PJ=0.0002 m=1 $X=75600 $Y=110300 $D=8
D140 DIO VDD_PAD dn PJ=0.0002 m=1 $X=77920 $Y=-95300 $D=8
D141 DIO VDD_PAD dn PJ=0.0002 m=1 $X=77920 $Y=114700 $D=8
D142 GND_PAD DIO dn PJ=0.0002 m=1 $X=80240 $Y=-99700 $D=8
D143 GND_PAD DIO dn PJ=0.0002 m=1 $X=80240 $Y=110300 $D=8
D144 DIO VDD_PAD dn PJ=0.0002 m=1 $X=82560 $Y=-95300 $D=8
D145 DIO VDD_PAD dn PJ=0.0002 m=1 $X=82560 $Y=114700 $D=8
D146 GND_PAD DIO dn PJ=0.0001 m=1 $X=84880 $Y=-99700 $D=8
D147 GND_PAD DIO dn PJ=0.0001 m=1 $X=84880 $Y=110300 $D=8
D148 DIO VDD_PAD dn PJ=0.0001 m=1 $X=88060 $Y=4700 $D=8
D149 DIO VDD_PAD dn PJ=0.0001 m=1 $X=88060 $Y=214700 $D=8
D150 GND_PAD DIO dn PJ=0.0002 m=1 $X=90380 $Y=-99700 $D=8
D151 GND_PAD DIO dn PJ=0.0002 m=1 $X=90380 $Y=110300 $D=8
D152 DIO VDD_PAD dn PJ=0.0002 m=1 $X=92700 $Y=-95300 $D=8
D153 DIO VDD_PAD dn PJ=0.0002 m=1 $X=92700 $Y=114700 $D=8
D154 GND_PAD DIO dn PJ=0.0002 m=1 $X=95020 $Y=-99700 $D=8
D155 GND_PAD DIO dn PJ=0.0002 m=1 $X=95020 $Y=110300 $D=8
D156 gnd! 36 dn PJ=5e-06 m=1 $X=1560 $Y=329900 $D=10
D157 36 vdd! dn PJ=5e-06 m=1 $X=1560 $Y=332220 $D=10
D158 gnd! 36 dn PJ=5e-06 m=1 $X=1560 $Y=328560 $D=11
D159 36 vdd! dn PJ=5e-06 m=1 $X=1560 $Y=334960 $D=11
X187 DIO 36 PAD $T=0 1440 0 0 $X=-5000 $Y=-235000
X188 27 28 34 pmos_a_CDNS_5887047866574 $T=78240 324220 0 0 $X=78240 $Y=324220
X189 vdd! 27 30 pmos_a_CDNS_5887047866574 $T=80480 324220 0 0 $X=80480 $Y=324220
X190 gnd! 11 28 nmos_a_CDNS_5887047866573 $T=75100 324160 0 0 $X=75100 $Y=324160
X191 gnd! 11 28 nmos_a_CDNS_5887047866573 $T=75100 331420 0 0 $X=75100 $Y=331420
X192 gnd! 26 29 nmos_a_CDNS_5887047866573 $T=77300 316840 0 0 $X=77300 $Y=316840
X193 gnd! 28 34 nmos_a_CDNS_5887047866573 $T=78240 330660 0 0 $X=78240 $Y=330660
X194 gnd! 28 30 nmos_a_CDNS_5887047866573 $T=80480 330660 0 0 $X=80480 $Y=330660
X195 gnd! 14 33 nmos_a_CDNS_5887047866586 $T=94080 316840 1 180 $X=91120 $Y=316840
X196 gnd! 12 33 nmos_a_CDNS_5887047866586 $T=94080 324400 1 180 $X=91120 $Y=324400
X199 vdd! 11 28 28 pmos_a_CDNS_5887047866592 $T=75100 323580 1 180 $X=71340 $Y=323580
X200 vdd! 11 28 28 pmos_a_CDNS_5887047866592 $T=75100 330880 1 180 $X=71340 $Y=330880
X201 vdd! 33 31 34 pmos_a_CDNS_5887047866592 $T=87320 332340 0 0 $X=87320 $Y=332340
X202 vdd! 12 33 33 pmos_a_CDNS_5887047866592 $T=87360 325000 0 0 $X=87360 $Y=325000
X203 GND_PAD DIO 12 nmos_io_a_CDNS_5887047866594 $T=13120 112700 0 0 $X=13120 $Y=112600
X204 GND_PAD DIO 12 nmos_io_a_CDNS_5887047866594 $T=13120 122340 0 0 $X=13120 $Y=122240
X205 GND_PAD DIO 12 nmos_io_a_CDNS_5887047866594 $T=13120 138700 0 0 $X=13120 $Y=138600
X206 GND_PAD DIO 12 nmos_io_a_CDNS_5887047866594 $T=13120 148340 0 0 $X=13120 $Y=148240
X207 GND_PAD DIO 12 nmos_io_a_CDNS_5887047866594 $T=13120 164700 0 0 $X=13120 $Y=164600
X208 GND_PAD DIO 12 nmos_io_a_CDNS_5887047866594 $T=13120 174340 0 0 $X=13120 $Y=174240
X209 GND_PAD DIO 12 nmos_io_a_CDNS_5887047866594 $T=13120 190700 0 0 $X=13120 $Y=190600
X210 GND_PAD DIO 12 nmos_io_a_CDNS_5887047866594 $T=13120 200340 0 0 $X=13120 $Y=200240
X211 GND_PAD DIO 12 nmos_io_a_CDNS_5887047866594 $T=27900 112700 0 0 $X=27900 $Y=112600
X212 GND_PAD DIO 12 nmos_io_a_CDNS_5887047866594 $T=27900 122340 0 0 $X=27900 $Y=122240
X213 GND_PAD DIO 12 nmos_io_a_CDNS_5887047866594 $T=27900 138700 0 0 $X=27900 $Y=138600
X214 GND_PAD DIO 12 nmos_io_a_CDNS_5887047866594 $T=27900 148340 0 0 $X=27900 $Y=148240
X215 GND_PAD DIO 12 nmos_io_a_CDNS_5887047866594 $T=27900 164700 0 0 $X=27900 $Y=164600
X216 GND_PAD DIO 12 nmos_io_a_CDNS_5887047866594 $T=27900 174340 0 0 $X=27900 $Y=174240
X217 GND_PAD DIO 12 nmos_io_a_CDNS_5887047866594 $T=27900 190700 0 0 $X=27900 $Y=190600
X218 GND_PAD DIO 12 nmos_io_a_CDNS_5887047866594 $T=27900 200340 0 0 $X=27900 $Y=200240
X219 GND_PAD DIO 12 nmos_io_a_CDNS_5887047866594 $T=42680 112700 0 0 $X=42680 $Y=112600
X220 GND_PAD DIO 12 nmos_io_a_CDNS_5887047866594 $T=42680 122340 0 0 $X=42680 $Y=122240
X221 GND_PAD DIO 12 nmos_io_a_CDNS_5887047866594 $T=42680 138700 0 0 $X=42680 $Y=138600
X222 GND_PAD DIO 12 nmos_io_a_CDNS_5887047866594 $T=42680 148340 0 0 $X=42680 $Y=148240
X223 GND_PAD DIO 12 nmos_io_a_CDNS_5887047866594 $T=42680 164700 0 0 $X=42680 $Y=164600
X224 GND_PAD DIO 12 nmos_io_a_CDNS_5887047866594 $T=42680 174340 0 0 $X=42680 $Y=174240
X225 GND_PAD DIO 12 nmos_io_a_CDNS_5887047866594 $T=42680 190700 0 0 $X=42680 $Y=190600
X226 GND_PAD DIO 12 nmos_io_a_CDNS_5887047866594 $T=42680 200340 0 0 $X=42680 $Y=200240
X227 GND_PAD DIO 14 nmos_io_a_CDNS_5887047866594 $T=57460 112700 0 0 $X=57460 $Y=112600
X228 GND_PAD DIO 14 nmos_io_a_CDNS_5887047866594 $T=57460 122340 0 0 $X=57460 $Y=122240
X229 GND_PAD DIO 14 nmos_io_a_CDNS_5887047866594 $T=57460 138700 0 0 $X=57460 $Y=138600
X230 GND_PAD DIO 14 nmos_io_a_CDNS_5887047866594 $T=57460 148340 0 0 $X=57460 $Y=148240
X231 GND_PAD DIO 14 nmos_io_a_CDNS_5887047866594 $T=57460 164700 0 0 $X=57460 $Y=164600
X232 GND_PAD DIO 14 nmos_io_a_CDNS_5887047866594 $T=57460 174340 0 0 $X=57460 $Y=174240
X233 GND_PAD DIO 14 nmos_io_a_CDNS_5887047866594 $T=57460 190700 0 0 $X=57460 $Y=190600
X234 GND_PAD DIO 14 nmos_io_a_CDNS_5887047866594 $T=57460 200340 0 0 $X=57460 $Y=200240
X235 GND_PAD DIO 14 nmos_io_a_CDNS_5887047866594 $T=72240 112700 0 0 $X=72240 $Y=112600
X236 GND_PAD DIO 14 nmos_io_a_CDNS_5887047866594 $T=72240 122340 0 0 $X=72240 $Y=122240
X237 GND_PAD DIO 14 nmos_io_a_CDNS_5887047866594 $T=72240 138700 0 0 $X=72240 $Y=138600
X238 GND_PAD DIO 14 nmos_io_a_CDNS_5887047866594 $T=72240 148340 0 0 $X=72240 $Y=148240
X239 GND_PAD DIO 14 nmos_io_a_CDNS_5887047866594 $T=72240 164700 0 0 $X=72240 $Y=164600
X240 GND_PAD DIO 14 nmos_io_a_CDNS_5887047866594 $T=72240 174340 0 0 $X=72240 $Y=174240
X241 GND_PAD DIO 14 nmos_io_a_CDNS_5887047866594 $T=72240 190700 0 0 $X=72240 $Y=190600
X242 GND_PAD DIO 14 nmos_io_a_CDNS_5887047866594 $T=72240 200340 0 0 $X=72240 $Y=200240
X243 GND_PAD DIO 14 nmos_io_a_CDNS_5887047866594 $T=87020 112700 0 0 $X=87020 $Y=112600
X244 GND_PAD DIO 14 nmos_io_a_CDNS_5887047866594 $T=87020 122340 0 0 $X=87020 $Y=122240
X245 GND_PAD DIO 14 nmos_io_a_CDNS_5887047866594 $T=87020 138700 0 0 $X=87020 $Y=138600
X246 GND_PAD DIO 14 nmos_io_a_CDNS_5887047866594 $T=87020 148340 0 0 $X=87020 $Y=148240
X247 GND_PAD DIO 14 nmos_io_a_CDNS_5887047866594 $T=87020 164700 0 0 $X=87020 $Y=164600
X248 GND_PAD DIO 14 nmos_io_a_CDNS_5887047866594 $T=87020 174340 0 0 $X=87020 $Y=174240
X249 GND_PAD DIO 14 nmos_io_a_CDNS_5887047866594 $T=87020 190700 0 0 $X=87020 $Y=190600
X250 GND_PAD DIO 14 nmos_io_a_CDNS_5887047866594 $T=87020 200340 0 0 $X=87020 $Y=200240
X251 29 gnd! dn_CDNS_5887047866588 $T=81960 318900 1 180 $X=80560 $Y=318600
X252 vdd! 29 dn_CDNS_5887047866588 $T=84440 318900 1 180 $X=83040 $Y=318600
X253 VDD_PAD DIO 11 pmos_io_a_CDNS_5887047866595 $T=13700 214500 1 180 $X=10800 $Y=214400
X254 VDD_PAD DIO 11 pmos_io_a_CDNS_5887047866595 $T=13700 226780 1 180 $X=10800 $Y=226680
X255 VDD_PAD DIO 11 pmos_io_a_CDNS_5887047866595 $T=13700 240500 1 180 $X=10800 $Y=240400
X256 VDD_PAD DIO 11 pmos_io_a_CDNS_5887047866595 $T=13700 252780 1 180 $X=10800 $Y=252680
X257 VDD_PAD DIO 11 pmos_io_a_CDNS_5887047866595 $T=13700 266500 1 180 $X=10800 $Y=266400
X258 VDD_PAD DIO 11 pmos_io_a_CDNS_5887047866595 $T=13700 278780 1 180 $X=10800 $Y=278680
X259 VDD_PAD DIO 11 pmos_io_a_CDNS_5887047866595 $T=13700 292500 1 180 $X=10800 $Y=292400
X260 VDD_PAD DIO 11 pmos_io_a_CDNS_5887047866595 $T=13700 304780 1 180 $X=10800 $Y=304680
X261 VDD_PAD DIO 11 pmos_io_a_CDNS_5887047866595 $T=28480 214500 1 180 $X=25580 $Y=214400
X262 VDD_PAD DIO 11 pmos_io_a_CDNS_5887047866595 $T=28480 226780 1 180 $X=25580 $Y=226680
X263 VDD_PAD DIO 11 pmos_io_a_CDNS_5887047866595 $T=28480 240500 1 180 $X=25580 $Y=240400
X264 VDD_PAD DIO 11 pmos_io_a_CDNS_5887047866595 $T=28480 252780 1 180 $X=25580 $Y=252680
X265 VDD_PAD DIO 11 pmos_io_a_CDNS_5887047866595 $T=28480 266500 1 180 $X=25580 $Y=266400
X266 VDD_PAD DIO 11 pmos_io_a_CDNS_5887047866595 $T=28480 278780 1 180 $X=25580 $Y=278680
X267 VDD_PAD DIO 11 pmos_io_a_CDNS_5887047866595 $T=28480 292500 1 180 $X=25580 $Y=292400
X268 VDD_PAD DIO 11 pmos_io_a_CDNS_5887047866595 $T=28480 304780 1 180 $X=25580 $Y=304680
X269 VDD_PAD DIO 11 pmos_io_a_CDNS_5887047866595 $T=43260 214500 1 180 $X=40360 $Y=214400
X270 VDD_PAD DIO 11 pmos_io_a_CDNS_5887047866595 $T=43260 226780 1 180 $X=40360 $Y=226680
X271 VDD_PAD DIO 11 pmos_io_a_CDNS_5887047866595 $T=43260 240500 1 180 $X=40360 $Y=240400
X272 VDD_PAD DIO 11 pmos_io_a_CDNS_5887047866595 $T=43260 252780 1 180 $X=40360 $Y=252680
X273 VDD_PAD DIO 11 pmos_io_a_CDNS_5887047866595 $T=43260 266500 1 180 $X=40360 $Y=266400
X274 VDD_PAD DIO 11 pmos_io_a_CDNS_5887047866595 $T=43260 278780 1 180 $X=40360 $Y=278680
X275 VDD_PAD DIO 11 pmos_io_a_CDNS_5887047866595 $T=43260 292500 1 180 $X=40360 $Y=292400
X276 VDD_PAD DIO 11 pmos_io_a_CDNS_5887047866595 $T=43260 304780 1 180 $X=40360 $Y=304680
X277 VDD_PAD DIO 13 pmos_io_a_CDNS_5887047866595 $T=58040 214500 1 180 $X=55140 $Y=214400
X278 VDD_PAD DIO 13 pmos_io_a_CDNS_5887047866595 $T=58040 226780 1 180 $X=55140 $Y=226680
X279 VDD_PAD DIO 13 pmos_io_a_CDNS_5887047866595 $T=58040 240500 1 180 $X=55140 $Y=240400
X280 VDD_PAD DIO 13 pmos_io_a_CDNS_5887047866595 $T=58040 252780 1 180 $X=55140 $Y=252680
X281 VDD_PAD DIO 13 pmos_io_a_CDNS_5887047866595 $T=58040 266500 1 180 $X=55140 $Y=266400
X282 VDD_PAD DIO 13 pmos_io_a_CDNS_5887047866595 $T=58040 278780 1 180 $X=55140 $Y=278680
X283 VDD_PAD DIO 13 pmos_io_a_CDNS_5887047866595 $T=58040 292500 1 180 $X=55140 $Y=292400
X284 VDD_PAD DIO 13 pmos_io_a_CDNS_5887047866595 $T=58040 304780 1 180 $X=55140 $Y=304680
X285 VDD_PAD DIO 13 pmos_io_a_CDNS_5887047866595 $T=72820 214500 1 180 $X=69920 $Y=214400
X286 VDD_PAD DIO 13 pmos_io_a_CDNS_5887047866595 $T=72820 226780 1 180 $X=69920 $Y=226680
X287 VDD_PAD DIO 13 pmos_io_a_CDNS_5887047866595 $T=72820 240500 1 180 $X=69920 $Y=240400
X288 VDD_PAD DIO 13 pmos_io_a_CDNS_5887047866595 $T=72820 252780 1 180 $X=69920 $Y=252680
X289 VDD_PAD DIO 13 pmos_io_a_CDNS_5887047866595 $T=72820 266500 1 180 $X=69920 $Y=266400
X290 VDD_PAD DIO 13 pmos_io_a_CDNS_5887047866595 $T=72820 278780 1 180 $X=69920 $Y=278680
X291 VDD_PAD DIO 13 pmos_io_a_CDNS_5887047866595 $T=72820 292500 1 180 $X=69920 $Y=292400
X292 VDD_PAD DIO 13 pmos_io_a_CDNS_5887047866595 $T=72820 304780 1 180 $X=69920 $Y=304680
X293 vdd! gnd! cpoly_n_CDNS_5887047866515 $T=16840 336500 0 0 $X=16840 $Y=336500
.ENDS
***************************************
.SUBCKT ICV_30 1 2 3 4 5 6 8 9 10
** N=10 EP=9 IP=14 FDC=2745
X0 1 2 3 4 PAD_Fill_200 $T=0 0 0 0 $X=0 $Y=-136000
X1 5 1 2 3 4 6 8 9 10 PADIO $T=0 100000 1 180 $X=-105000 $Y=-135000
.ENDS
***************************************
.SUBCKT dn_CDNS_588704786652
** N=2 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT ICV_31 1 2 3
** N=3 EP=3 IP=4 FDC=2
D0 2 3 dn PJ=0.00041 m=1 $X=2740 $Y=0 $D=8
D1 2 1 dn PJ=0.00041 m=1 $X=-460 $Y=0 $D=9
.ENDS
***************************************
.SUBCKT ICV_32 1 2
** N=2 EP=2 IP=6 FDC=4
X0 1 2 1 ICV_31 $T=0 0 0 0 $X=-640 $Y=-300
X1 1 2 1 ICV_31 $T=5000 0 0 0 $X=4360 $Y=-300
.ENDS
***************************************
.SUBCKT ICV_33 1 2
** N=2 EP=2 IP=4 FDC=8
X0 1 2 ICV_32 $T=0 0 0 0 $X=-640 $Y=-300
X1 1 2 ICV_32 $T=10000 0 0 0 $X=9360 $Y=-300
.ENDS
***************************************
.SUBCKT GND_Core gnd vdd!
** N=6 EP=2 IP=16 FDC=115
D0 gnd vdd! dn PJ=0.00041 m=1 $X=94280 $Y=-99700 $D=9
X1 vdd! gnd cpoly_n_CDNS_588704786651 $T=520 333340 0 0 $X=520 $Y=333340
X2 gnd vdd! cpoly_p_CDNS_588704786650 $T=520 320500 0 0 $X=520 $Y=320500
X4 vdd! gnd ICV_32 $T=84740 -99700 0 0 $X=84100 $Y=-100000
X5 vdd! gnd ICV_33 $T=4740 -99700 0 0 $X=4100 $Y=-100000
X6 vdd! gnd ICV_33 $T=24740 -99700 0 0 $X=24100 $Y=-100000
X7 vdd! gnd ICV_33 $T=44740 -99700 0 0 $X=44100 $Y=-100000
X8 vdd! gnd ICV_33 $T=64740 -99700 0 0 $X=64100 $Y=-100000
.ENDS
***************************************
.SUBCKT nmos_io_a_CDNS_5887047866531 1 2 3
** N=3 EP=3 IP=0 FDC=1
M0 2 3 1 1 nmos_io_a L=2.8e-07 W=1e-05 AD=7.39066e-12 AS=2.5056e-13 PD=4.0608e-06 PS=2.0304e-06 w_cont=4.1e-06 nfing=1 $X=620 $Y=200 $D=0
.ENDS
***************************************
.SUBCKT cpoly_n_CDNS_5887047866535 1 2
** N=2 EP=2 IP=0 FDC=80
M0 1 2 1 cpoly_n w=6e-06 l=2e-06 c=7.5402e-14 as=2.4e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.4338e-06 sim_w=5.76e-06 m_per_maxw=1.04167 numb_sub_cont=3 nfing=1 $X=620 $Y=200 $D=22
M1 1 2 1 cpoly_n w=6e-06 l=2e-06 c=7.5402e-14 as=3.0336e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.4338e-06 sim_w=5.76e-06 m_per_maxw=1.04167 numb_sub_cont=3 nfing=1 $X=3140 $Y=200 $D=22
M2 1 2 1 cpoly_n w=6e-06 l=2e-06 c=7.5402e-14 as=3.0336e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.4338e-06 sim_w=5.76e-06 m_per_maxw=1.04167 numb_sub_cont=3 nfing=1 $X=5660 $Y=200 $D=22
M3 1 2 1 cpoly_n w=6e-06 l=2e-06 c=7.5402e-14 as=3.0336e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.4338e-06 sim_w=5.76e-06 m_per_maxw=1.04167 numb_sub_cont=3 nfing=1 $X=8180 $Y=200 $D=22
M4 1 2 1 cpoly_n w=6e-06 l=2e-06 c=7.5402e-14 as=3.0336e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.4338e-06 sim_w=5.76e-06 m_per_maxw=1.04167 numb_sub_cont=3 nfing=1 $X=10700 $Y=200 $D=22
M5 1 2 1 cpoly_n w=6e-06 l=2e-06 c=7.5402e-14 as=3.0336e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.4338e-06 sim_w=5.76e-06 m_per_maxw=1.04167 numb_sub_cont=3 nfing=1 $X=13220 $Y=200 $D=22
M6 1 2 1 cpoly_n w=6e-06 l=2e-06 c=7.5402e-14 as=3.0336e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.4338e-06 sim_w=5.76e-06 m_per_maxw=1.04167 numb_sub_cont=3 nfing=1 $X=15740 $Y=200 $D=22
M7 1 2 1 cpoly_n w=6e-06 l=2e-06 c=7.5402e-14 as=3.0336e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.4338e-06 sim_w=5.76e-06 m_per_maxw=1.04167 numb_sub_cont=3 nfing=1 $X=18260 $Y=200 $D=22
M8 1 2 1 cpoly_n w=6e-06 l=2e-06 c=7.5402e-14 as=3.0336e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.4338e-06 sim_w=5.76e-06 m_per_maxw=1.04167 numb_sub_cont=3 nfing=1 $X=20780 $Y=200 $D=22
M9 1 2 1 cpoly_n w=6e-06 l=2e-06 c=7.5402e-14 as=3.0336e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.4338e-06 sim_w=5.76e-06 m_per_maxw=1.04167 numb_sub_cont=3 nfing=1 $X=23300 $Y=200 $D=22
M10 1 2 1 cpoly_n w=6e-06 l=2e-06 c=7.5402e-14 as=3.0336e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.4338e-06 sim_w=5.76e-06 m_per_maxw=1.04167 numb_sub_cont=3 nfing=1 $X=25820 $Y=200 $D=22
M11 1 2 1 cpoly_n w=6e-06 l=2e-06 c=7.5402e-14 as=3.0336e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.4338e-06 sim_w=5.76e-06 m_per_maxw=1.04167 numb_sub_cont=3 nfing=1 $X=28340 $Y=200 $D=22
M12 1 2 1 cpoly_n w=6e-06 l=2e-06 c=7.5402e-14 as=3.0336e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.4338e-06 sim_w=5.76e-06 m_per_maxw=1.04167 numb_sub_cont=3 nfing=1 $X=30860 $Y=200 $D=22
M13 1 2 1 cpoly_n w=6e-06 l=2e-06 c=7.5402e-14 as=3.0336e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.4338e-06 sim_w=5.76e-06 m_per_maxw=1.04167 numb_sub_cont=3 nfing=1 $X=33380 $Y=200 $D=22
M14 1 2 1 cpoly_n w=6e-06 l=2e-06 c=7.5402e-14 as=3.0336e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.4338e-06 sim_w=5.76e-06 m_per_maxw=1.04167 numb_sub_cont=3 nfing=1 $X=35900 $Y=200 $D=22
M15 1 2 1 cpoly_n w=6e-06 l=2e-06 c=7.5402e-14 as=3.0336e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.4338e-06 sim_w=5.76e-06 m_per_maxw=1.04167 numb_sub_cont=3 nfing=1 $X=38420 $Y=200 $D=22
M16 1 2 1 cpoly_n w=6e-06 l=2e-06 c=7.5402e-14 as=3.0336e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.4338e-06 sim_w=5.76e-06 m_per_maxw=1.04167 numb_sub_cont=3 nfing=1 $X=40940 $Y=200 $D=22
M17 1 2 1 cpoly_n w=6e-06 l=2e-06 c=7.5402e-14 as=3.0336e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.4338e-06 sim_w=5.76e-06 m_per_maxw=1.04167 numb_sub_cont=3 nfing=1 $X=43460 $Y=200 $D=22
M18 1 2 1 cpoly_n w=6e-06 l=2e-06 c=7.5402e-14 as=3.0336e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.4338e-06 sim_w=5.76e-06 m_per_maxw=1.04167 numb_sub_cont=3 nfing=1 $X=45980 $Y=200 $D=22
M19 1 2 1 cpoly_n w=6e-06 l=2e-06 c=7.5402e-14 as=3.0336e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.4338e-06 sim_w=5.76e-06 m_per_maxw=1.04167 numb_sub_cont=3 nfing=1 $X=48500 $Y=200 $D=22
M20 1 2 1 cpoly_n w=6e-06 l=2e-06 c=7.5402e-14 as=3.0336e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.4338e-06 sim_w=5.76e-06 m_per_maxw=1.04167 numb_sub_cont=3 nfing=1 $X=51020 $Y=200 $D=22
M21 1 2 1 cpoly_n w=6e-06 l=2e-06 c=7.5402e-14 as=3.0336e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.4338e-06 sim_w=5.76e-06 m_per_maxw=1.04167 numb_sub_cont=3 nfing=1 $X=53540 $Y=200 $D=22
M22 1 2 1 cpoly_n w=6e-06 l=2e-06 c=7.5402e-14 as=3.0336e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.4338e-06 sim_w=5.76e-06 m_per_maxw=1.04167 numb_sub_cont=3 nfing=1 $X=56060 $Y=200 $D=22
M23 1 2 1 cpoly_n w=6e-06 l=2e-06 c=7.5402e-14 as=3.0336e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.4338e-06 sim_w=5.76e-06 m_per_maxw=1.04167 numb_sub_cont=3 nfing=1 $X=58580 $Y=200 $D=22
M24 1 2 1 cpoly_n w=6e-06 l=2e-06 c=7.5402e-14 as=3.0336e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.4338e-06 sim_w=5.76e-06 m_per_maxw=1.04167 numb_sub_cont=3 nfing=1 $X=61100 $Y=200 $D=22
M25 1 2 1 cpoly_n w=6e-06 l=2e-06 c=7.5402e-14 as=3.0336e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.4338e-06 sim_w=5.76e-06 m_per_maxw=1.04167 numb_sub_cont=3 nfing=1 $X=63620 $Y=200 $D=22
M26 1 2 1 cpoly_n w=6e-06 l=2e-06 c=7.5402e-14 as=3.0336e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.4338e-06 sim_w=5.76e-06 m_per_maxw=1.04167 numb_sub_cont=3 nfing=1 $X=66140 $Y=200 $D=22
M27 1 2 1 cpoly_n w=6e-06 l=2e-06 c=7.5402e-14 as=3.0336e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.4338e-06 sim_w=5.76e-06 m_per_maxw=1.04167 numb_sub_cont=3 nfing=1 $X=68660 $Y=200 $D=22
M28 1 2 1 cpoly_n w=6e-06 l=2e-06 c=7.5402e-14 as=3.0336e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.4338e-06 sim_w=5.76e-06 m_per_maxw=1.04167 numb_sub_cont=3 nfing=1 $X=71180 $Y=200 $D=22
M29 1 2 1 cpoly_n w=6e-06 l=2e-06 c=7.5402e-14 as=3.0336e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.4338e-06 sim_w=5.76e-06 m_per_maxw=1.04167 numb_sub_cont=3 nfing=1 $X=73700 $Y=200 $D=22
M30 1 2 1 cpoly_n w=6e-06 l=2e-06 c=7.5402e-14 as=3.0336e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.4338e-06 sim_w=5.76e-06 m_per_maxw=1.04167 numb_sub_cont=3 nfing=1 $X=76220 $Y=200 $D=22
M31 1 2 1 cpoly_n w=6e-06 l=2e-06 c=7.5402e-14 as=3.0336e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.4338e-06 sim_w=5.76e-06 m_per_maxw=1.04167 numb_sub_cont=3 nfing=1 $X=78740 $Y=200 $D=22
M32 1 2 1 cpoly_n w=6e-06 l=2e-06 c=7.5402e-14 as=3.0336e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.4338e-06 sim_w=5.76e-06 m_per_maxw=1.04167 numb_sub_cont=3 nfing=1 $X=81260 $Y=200 $D=22
M33 1 2 1 cpoly_n w=6e-06 l=2e-06 c=7.5402e-14 as=3.0336e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.4338e-06 sim_w=5.76e-06 m_per_maxw=1.04167 numb_sub_cont=3 nfing=1 $X=83780 $Y=200 $D=22
M34 1 2 1 cpoly_n w=6e-06 l=2e-06 c=7.5402e-14 as=3.0336e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.4338e-06 sim_w=5.76e-06 m_per_maxw=1.04167 numb_sub_cont=3 nfing=1 $X=86300 $Y=200 $D=22
M35 1 2 1 cpoly_n w=6e-06 l=2e-06 c=7.5402e-14 as=3.0336e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.4338e-06 sim_w=5.76e-06 m_per_maxw=1.04167 numb_sub_cont=3 nfing=1 $X=88820 $Y=200 $D=22
M36 1 2 1 cpoly_n w=6e-06 l=2e-06 c=7.5402e-14 as=3.0336e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.4338e-06 sim_w=5.76e-06 m_per_maxw=1.04167 numb_sub_cont=3 nfing=1 $X=91340 $Y=200 $D=22
M37 1 2 1 cpoly_n w=6e-06 l=2e-06 c=7.5402e-14 as=3.0336e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.4338e-06 sim_w=5.76e-06 m_per_maxw=1.04167 numb_sub_cont=3 nfing=1 $X=93860 $Y=200 $D=22
M38 1 2 1 cpoly_n w=6e-06 l=2e-06 c=7.5402e-14 as=3.0336e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.4338e-06 sim_w=5.76e-06 m_per_maxw=1.04167 numb_sub_cont=3 nfing=1 $X=96380 $Y=200 $D=22
M39 1 2 1 cpoly_n w=6e-06 l=2e-06 c=7.5402e-14 as=3.0336e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.4338e-06 sim_w=5.76e-06 m_per_maxw=1.04167 numb_sub_cont=3 nfing=1 $X=98900 $Y=200 $D=22
M40 1 2 1 cpoly_n w=6e-06 l=2e-06 c=7.5402e-14 as=3.0336e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.4338e-06 sim_w=5.76e-06 m_per_maxw=1.04167 numb_sub_cont=3 nfing=1 $X=101420 $Y=200 $D=22
M41 1 2 1 cpoly_n w=6e-06 l=2e-06 c=7.5402e-14 as=3.0336e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.4338e-06 sim_w=5.76e-06 m_per_maxw=1.04167 numb_sub_cont=3 nfing=1 $X=103940 $Y=200 $D=22
M42 1 2 1 cpoly_n w=6e-06 l=2e-06 c=7.5402e-14 as=3.0336e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.4338e-06 sim_w=5.76e-06 m_per_maxw=1.04167 numb_sub_cont=3 nfing=1 $X=106460 $Y=200 $D=22
M43 1 2 1 cpoly_n w=6e-06 l=2e-06 c=7.5402e-14 as=3.0336e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.4338e-06 sim_w=5.76e-06 m_per_maxw=1.04167 numb_sub_cont=3 nfing=1 $X=108980 $Y=200 $D=22
M44 1 2 1 cpoly_n w=6e-06 l=2e-06 c=7.5402e-14 as=3.0336e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.4338e-06 sim_w=5.76e-06 m_per_maxw=1.04167 numb_sub_cont=3 nfing=1 $X=111500 $Y=200 $D=22
M45 1 2 1 cpoly_n w=6e-06 l=2e-06 c=7.5402e-14 as=3.0336e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.4338e-06 sim_w=5.76e-06 m_per_maxw=1.04167 numb_sub_cont=3 nfing=1 $X=114020 $Y=200 $D=22
M46 1 2 1 cpoly_n w=6e-06 l=2e-06 c=7.5402e-14 as=3.0336e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.4338e-06 sim_w=5.76e-06 m_per_maxw=1.04167 numb_sub_cont=3 nfing=1 $X=116540 $Y=200 $D=22
M47 1 2 1 cpoly_n w=6e-06 l=2e-06 c=7.5402e-14 as=3.0336e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.4338e-06 sim_w=5.76e-06 m_per_maxw=1.04167 numb_sub_cont=3 nfing=1 $X=119060 $Y=200 $D=22
M48 1 2 1 cpoly_n w=6e-06 l=2e-06 c=7.5402e-14 as=3.0336e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.4338e-06 sim_w=5.76e-06 m_per_maxw=1.04167 numb_sub_cont=3 nfing=1 $X=121580 $Y=200 $D=22
M49 1 2 1 cpoly_n w=6e-06 l=2e-06 c=7.5402e-14 as=3.0336e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.4338e-06 sim_w=5.76e-06 m_per_maxw=1.04167 numb_sub_cont=3 nfing=1 $X=124100 $Y=200 $D=22
M50 1 2 1 cpoly_n w=6e-06 l=2e-06 c=7.5402e-14 as=3.0336e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.4338e-06 sim_w=5.76e-06 m_per_maxw=1.04167 numb_sub_cont=3 nfing=1 $X=126620 $Y=200 $D=22
M51 1 2 1 cpoly_n w=6e-06 l=2e-06 c=7.5402e-14 as=3.0336e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.4338e-06 sim_w=5.76e-06 m_per_maxw=1.04167 numb_sub_cont=3 nfing=1 $X=129140 $Y=200 $D=22
M52 1 2 1 cpoly_n w=6e-06 l=2e-06 c=7.5402e-14 as=3.0336e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.4338e-06 sim_w=5.76e-06 m_per_maxw=1.04167 numb_sub_cont=3 nfing=1 $X=131660 $Y=200 $D=22
M53 1 2 1 cpoly_n w=6e-06 l=2e-06 c=7.5402e-14 as=3.0336e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.4338e-06 sim_w=5.76e-06 m_per_maxw=1.04167 numb_sub_cont=3 nfing=1 $X=134180 $Y=200 $D=22
M54 1 2 1 cpoly_n w=6e-06 l=2e-06 c=7.5402e-14 as=3.0336e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.4338e-06 sim_w=5.76e-06 m_per_maxw=1.04167 numb_sub_cont=3 nfing=1 $X=136700 $Y=200 $D=22
M55 1 2 1 cpoly_n w=6e-06 l=2e-06 c=7.5402e-14 as=3.0336e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.4338e-06 sim_w=5.76e-06 m_per_maxw=1.04167 numb_sub_cont=3 nfing=1 $X=139220 $Y=200 $D=22
M56 1 2 1 cpoly_n w=6e-06 l=2e-06 c=7.5402e-14 as=3.0336e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.4338e-06 sim_w=5.76e-06 m_per_maxw=1.04167 numb_sub_cont=3 nfing=1 $X=141740 $Y=200 $D=22
M57 1 2 1 cpoly_n w=6e-06 l=2e-06 c=7.5402e-14 as=3.0336e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.4338e-06 sim_w=5.76e-06 m_per_maxw=1.04167 numb_sub_cont=3 nfing=1 $X=144260 $Y=200 $D=22
M58 1 2 1 cpoly_n w=6e-06 l=2e-06 c=7.5402e-14 as=3.0336e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.4338e-06 sim_w=5.76e-06 m_per_maxw=1.04167 numb_sub_cont=3 nfing=1 $X=146780 $Y=200 $D=22
M59 1 2 1 cpoly_n w=6e-06 l=2e-06 c=7.5402e-14 as=3.0336e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.4338e-06 sim_w=5.76e-06 m_per_maxw=1.04167 numb_sub_cont=3 nfing=1 $X=149300 $Y=200 $D=22
M60 1 2 1 cpoly_n w=6e-06 l=2e-06 c=7.5402e-14 as=3.0336e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.4338e-06 sim_w=5.76e-06 m_per_maxw=1.04167 numb_sub_cont=3 nfing=1 $X=151820 $Y=200 $D=22
M61 1 2 1 cpoly_n w=6e-06 l=2e-06 c=7.5402e-14 as=3.0336e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.4338e-06 sim_w=5.76e-06 m_per_maxw=1.04167 numb_sub_cont=3 nfing=1 $X=154340 $Y=200 $D=22
M62 1 2 1 cpoly_n w=6e-06 l=2e-06 c=7.5402e-14 as=3.0336e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.4338e-06 sim_w=5.76e-06 m_per_maxw=1.04167 numb_sub_cont=3 nfing=1 $X=156860 $Y=200 $D=22
M63 1 2 1 cpoly_n w=6e-06 l=2e-06 c=7.5402e-14 as=3.0336e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.4338e-06 sim_w=5.76e-06 m_per_maxw=1.04167 numb_sub_cont=3 nfing=1 $X=159380 $Y=200 $D=22
M64 1 2 1 cpoly_n w=6e-06 l=2e-06 c=7.5402e-14 as=3.0336e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.4338e-06 sim_w=5.76e-06 m_per_maxw=1.04167 numb_sub_cont=3 nfing=1 $X=161900 $Y=200 $D=22
M65 1 2 1 cpoly_n w=6e-06 l=2e-06 c=7.5402e-14 as=3.0336e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.4338e-06 sim_w=5.76e-06 m_per_maxw=1.04167 numb_sub_cont=3 nfing=1 $X=164420 $Y=200 $D=22
M66 1 2 1 cpoly_n w=6e-06 l=2e-06 c=7.5402e-14 as=3.0336e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.4338e-06 sim_w=5.76e-06 m_per_maxw=1.04167 numb_sub_cont=3 nfing=1 $X=166940 $Y=200 $D=22
M67 1 2 1 cpoly_n w=6e-06 l=2e-06 c=7.5402e-14 as=3.0336e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.4338e-06 sim_w=5.76e-06 m_per_maxw=1.04167 numb_sub_cont=3 nfing=1 $X=169460 $Y=200 $D=22
M68 1 2 1 cpoly_n w=6e-06 l=2e-06 c=7.5402e-14 as=3.0336e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.4338e-06 sim_w=5.76e-06 m_per_maxw=1.04167 numb_sub_cont=3 nfing=1 $X=171980 $Y=200 $D=22
M69 1 2 1 cpoly_n w=6e-06 l=2e-06 c=7.5402e-14 as=3.0336e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.4338e-06 sim_w=5.76e-06 m_per_maxw=1.04167 numb_sub_cont=3 nfing=1 $X=174500 $Y=200 $D=22
M70 1 2 1 cpoly_n w=6e-06 l=2e-06 c=7.5402e-14 as=3.0336e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.4338e-06 sim_w=5.76e-06 m_per_maxw=1.04167 numb_sub_cont=3 nfing=1 $X=177020 $Y=200 $D=22
M71 1 2 1 cpoly_n w=6e-06 l=2e-06 c=7.5402e-14 as=3.0336e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.4338e-06 sim_w=5.76e-06 m_per_maxw=1.04167 numb_sub_cont=3 nfing=1 $X=179540 $Y=200 $D=22
M72 1 2 1 cpoly_n w=6e-06 l=2e-06 c=7.5402e-14 as=3.0336e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.4338e-06 sim_w=5.76e-06 m_per_maxw=1.04167 numb_sub_cont=3 nfing=1 $X=182060 $Y=200 $D=22
M73 1 2 1 cpoly_n w=6e-06 l=2e-06 c=7.5402e-14 as=3.0336e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.4338e-06 sim_w=5.76e-06 m_per_maxw=1.04167 numb_sub_cont=3 nfing=1 $X=184580 $Y=200 $D=22
M74 1 2 1 cpoly_n w=6e-06 l=2e-06 c=7.5402e-14 as=3.0336e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.4338e-06 sim_w=5.76e-06 m_per_maxw=1.04167 numb_sub_cont=3 nfing=1 $X=187100 $Y=200 $D=22
M75 1 2 1 cpoly_n w=6e-06 l=2e-06 c=7.5402e-14 as=3.0336e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.4338e-06 sim_w=5.76e-06 m_per_maxw=1.04167 numb_sub_cont=3 nfing=1 $X=189620 $Y=200 $D=22
M76 1 2 1 cpoly_n w=6e-06 l=2e-06 c=7.5402e-14 as=3.0336e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.4338e-06 sim_w=5.76e-06 m_per_maxw=1.04167 numb_sub_cont=3 nfing=1 $X=192140 $Y=200 $D=22
M77 1 2 1 cpoly_n w=6e-06 l=2e-06 c=7.5402e-14 as=3.0336e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.4338e-06 sim_w=5.76e-06 m_per_maxw=1.04167 numb_sub_cont=3 nfing=1 $X=194660 $Y=200 $D=22
M78 1 2 1 cpoly_n w=6e-06 l=2e-06 c=7.5402e-14 as=3.0336e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.4338e-06 sim_w=5.76e-06 m_per_maxw=1.04167 numb_sub_cont=3 nfing=1 $X=197180 $Y=200 $D=22
M79 1 2 1 cpoly_n w=6e-06 l=2e-06 c=7.5402e-14 as=2.4e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.4338e-06 sim_w=5.76e-06 m_per_maxw=1.04167 numb_sub_cont=3 nfing=1 $X=199700 $Y=200 $D=22
.ENDS
***************************************
.SUBCKT nmos_a_CDNS_5887047866530 1 2 3
** N=3 EP=3 IP=0 FDC=1
M0 2 3 1 1 nmos_a L=2.4e-07 W=4e-06 AD=1.7568e-12 AS=1.6e-12 PD=4.392e-06 PS=2.196e-06 w_cont=2.1e-06 nfing=1 source_num=2 $X=620 $Y=200 $D=1
.ENDS
***************************************
.SUBCKT cpoly_p_CDNS_5887047866528 1 2
** N=2 EP=2 IP=0 FDC=80
M0 1 2 1 cpoly_p w=6e-06 l=2e-06 c=8.0712e-14 as=1.68e-13 ad=7.488e-13 ps=1.44e-06 pd=1.13684e-06 sim_w=2.88e-06 m_per_maxw=2.08333 numb_sub_cont=4 nfing=1 $X=620 $Y=200 $D=21
M1 1 2 1 cpoly_p w=6e-06 l=2e-06 c=8.0712e-14 as=2.1408e-13 ad=7.488e-13 ps=1.44e-06 pd=1.13684e-06 sim_w=2.88e-06 m_per_maxw=2.08333 numb_sub_cont=4 nfing=1 $X=3140 $Y=200 $D=21
M2 1 2 1 cpoly_p w=6e-06 l=2e-06 c=8.0712e-14 as=2.1408e-13 ad=7.488e-13 ps=1.44e-06 pd=1.13684e-06 sim_w=2.88e-06 m_per_maxw=2.08333 numb_sub_cont=4 nfing=1 $X=5660 $Y=200 $D=21
M3 1 2 1 cpoly_p w=6e-06 l=2e-06 c=8.0712e-14 as=2.1408e-13 ad=7.488e-13 ps=1.44e-06 pd=1.13684e-06 sim_w=2.88e-06 m_per_maxw=2.08333 numb_sub_cont=4 nfing=1 $X=8180 $Y=200 $D=21
M4 1 2 1 cpoly_p w=6e-06 l=2e-06 c=8.0712e-14 as=2.1408e-13 ad=7.488e-13 ps=1.44e-06 pd=1.13684e-06 sim_w=2.88e-06 m_per_maxw=2.08333 numb_sub_cont=4 nfing=1 $X=10700 $Y=200 $D=21
M5 1 2 1 cpoly_p w=6e-06 l=2e-06 c=8.0712e-14 as=2.1408e-13 ad=7.488e-13 ps=1.44e-06 pd=1.13684e-06 sim_w=2.88e-06 m_per_maxw=2.08333 numb_sub_cont=4 nfing=1 $X=13220 $Y=200 $D=21
M6 1 2 1 cpoly_p w=6e-06 l=2e-06 c=8.0712e-14 as=2.1408e-13 ad=7.488e-13 ps=1.44e-06 pd=1.13684e-06 sim_w=2.88e-06 m_per_maxw=2.08333 numb_sub_cont=4 nfing=1 $X=15740 $Y=200 $D=21
M7 1 2 1 cpoly_p w=6e-06 l=2e-06 c=8.0712e-14 as=2.1408e-13 ad=7.488e-13 ps=1.44e-06 pd=1.13684e-06 sim_w=2.88e-06 m_per_maxw=2.08333 numb_sub_cont=4 nfing=1 $X=18260 $Y=200 $D=21
M8 1 2 1 cpoly_p w=6e-06 l=2e-06 c=8.0712e-14 as=2.1408e-13 ad=7.488e-13 ps=1.44e-06 pd=1.13684e-06 sim_w=2.88e-06 m_per_maxw=2.08333 numb_sub_cont=4 nfing=1 $X=20780 $Y=200 $D=21
M9 1 2 1 cpoly_p w=6e-06 l=2e-06 c=8.0712e-14 as=2.1408e-13 ad=7.488e-13 ps=1.44e-06 pd=1.13684e-06 sim_w=2.88e-06 m_per_maxw=2.08333 numb_sub_cont=4 nfing=1 $X=23300 $Y=200 $D=21
M10 1 2 1 cpoly_p w=6e-06 l=2e-06 c=8.0712e-14 as=2.1408e-13 ad=7.488e-13 ps=1.44e-06 pd=1.13684e-06 sim_w=2.88e-06 m_per_maxw=2.08333 numb_sub_cont=4 nfing=1 $X=25820 $Y=200 $D=21
M11 1 2 1 cpoly_p w=6e-06 l=2e-06 c=8.0712e-14 as=2.1408e-13 ad=7.488e-13 ps=1.44e-06 pd=1.13684e-06 sim_w=2.88e-06 m_per_maxw=2.08333 numb_sub_cont=4 nfing=1 $X=28340 $Y=200 $D=21
M12 1 2 1 cpoly_p w=6e-06 l=2e-06 c=8.0712e-14 as=2.1408e-13 ad=7.488e-13 ps=1.44e-06 pd=1.13684e-06 sim_w=2.88e-06 m_per_maxw=2.08333 numb_sub_cont=4 nfing=1 $X=30860 $Y=200 $D=21
M13 1 2 1 cpoly_p w=6e-06 l=2e-06 c=8.0712e-14 as=2.1408e-13 ad=7.488e-13 ps=1.44e-06 pd=1.13684e-06 sim_w=2.88e-06 m_per_maxw=2.08333 numb_sub_cont=4 nfing=1 $X=33380 $Y=200 $D=21
M14 1 2 1 cpoly_p w=6e-06 l=2e-06 c=8.0712e-14 as=2.1408e-13 ad=7.488e-13 ps=1.44e-06 pd=1.13684e-06 sim_w=2.88e-06 m_per_maxw=2.08333 numb_sub_cont=4 nfing=1 $X=35900 $Y=200 $D=21
M15 1 2 1 cpoly_p w=6e-06 l=2e-06 c=8.0712e-14 as=2.1408e-13 ad=7.488e-13 ps=1.44e-06 pd=1.13684e-06 sim_w=2.88e-06 m_per_maxw=2.08333 numb_sub_cont=4 nfing=1 $X=38420 $Y=200 $D=21
M16 1 2 1 cpoly_p w=6e-06 l=2e-06 c=8.0712e-14 as=2.1408e-13 ad=7.488e-13 ps=1.44e-06 pd=1.13684e-06 sim_w=2.88e-06 m_per_maxw=2.08333 numb_sub_cont=4 nfing=1 $X=40940 $Y=200 $D=21
M17 1 2 1 cpoly_p w=6e-06 l=2e-06 c=8.0712e-14 as=2.1408e-13 ad=7.488e-13 ps=1.44e-06 pd=1.13684e-06 sim_w=2.88e-06 m_per_maxw=2.08333 numb_sub_cont=4 nfing=1 $X=43460 $Y=200 $D=21
M18 1 2 1 cpoly_p w=6e-06 l=2e-06 c=8.0712e-14 as=2.1408e-13 ad=7.488e-13 ps=1.44e-06 pd=1.13684e-06 sim_w=2.88e-06 m_per_maxw=2.08333 numb_sub_cont=4 nfing=1 $X=45980 $Y=200 $D=21
M19 1 2 1 cpoly_p w=6e-06 l=2e-06 c=8.0712e-14 as=2.1408e-13 ad=7.488e-13 ps=1.44e-06 pd=1.13684e-06 sim_w=2.88e-06 m_per_maxw=2.08333 numb_sub_cont=4 nfing=1 $X=48500 $Y=200 $D=21
M20 1 2 1 cpoly_p w=6e-06 l=2e-06 c=8.0712e-14 as=2.1408e-13 ad=7.488e-13 ps=1.44e-06 pd=1.13684e-06 sim_w=2.88e-06 m_per_maxw=2.08333 numb_sub_cont=4 nfing=1 $X=51020 $Y=200 $D=21
M21 1 2 1 cpoly_p w=6e-06 l=2e-06 c=8.0712e-14 as=2.1408e-13 ad=7.488e-13 ps=1.44e-06 pd=1.13684e-06 sim_w=2.88e-06 m_per_maxw=2.08333 numb_sub_cont=4 nfing=1 $X=53540 $Y=200 $D=21
M22 1 2 1 cpoly_p w=6e-06 l=2e-06 c=8.0712e-14 as=2.1408e-13 ad=7.488e-13 ps=1.44e-06 pd=1.13684e-06 sim_w=2.88e-06 m_per_maxw=2.08333 numb_sub_cont=4 nfing=1 $X=56060 $Y=200 $D=21
M23 1 2 1 cpoly_p w=6e-06 l=2e-06 c=8.0712e-14 as=2.1408e-13 ad=7.488e-13 ps=1.44e-06 pd=1.13684e-06 sim_w=2.88e-06 m_per_maxw=2.08333 numb_sub_cont=4 nfing=1 $X=58580 $Y=200 $D=21
M24 1 2 1 cpoly_p w=6e-06 l=2e-06 c=8.0712e-14 as=2.1408e-13 ad=7.488e-13 ps=1.44e-06 pd=1.13684e-06 sim_w=2.88e-06 m_per_maxw=2.08333 numb_sub_cont=4 nfing=1 $X=61100 $Y=200 $D=21
M25 1 2 1 cpoly_p w=6e-06 l=2e-06 c=8.0712e-14 as=2.1408e-13 ad=7.488e-13 ps=1.44e-06 pd=1.13684e-06 sim_w=2.88e-06 m_per_maxw=2.08333 numb_sub_cont=4 nfing=1 $X=63620 $Y=200 $D=21
M26 1 2 1 cpoly_p w=6e-06 l=2e-06 c=8.0712e-14 as=2.1408e-13 ad=7.488e-13 ps=1.44e-06 pd=1.13684e-06 sim_w=2.88e-06 m_per_maxw=2.08333 numb_sub_cont=4 nfing=1 $X=66140 $Y=200 $D=21
M27 1 2 1 cpoly_p w=6e-06 l=2e-06 c=8.0712e-14 as=2.1408e-13 ad=7.488e-13 ps=1.44e-06 pd=1.13684e-06 sim_w=2.88e-06 m_per_maxw=2.08333 numb_sub_cont=4 nfing=1 $X=68660 $Y=200 $D=21
M28 1 2 1 cpoly_p w=6e-06 l=2e-06 c=8.0712e-14 as=2.1408e-13 ad=7.488e-13 ps=1.44e-06 pd=1.13684e-06 sim_w=2.88e-06 m_per_maxw=2.08333 numb_sub_cont=4 nfing=1 $X=71180 $Y=200 $D=21
M29 1 2 1 cpoly_p w=6e-06 l=2e-06 c=8.0712e-14 as=2.1408e-13 ad=7.488e-13 ps=1.44e-06 pd=1.13684e-06 sim_w=2.88e-06 m_per_maxw=2.08333 numb_sub_cont=4 nfing=1 $X=73700 $Y=200 $D=21
M30 1 2 1 cpoly_p w=6e-06 l=2e-06 c=8.0712e-14 as=2.1408e-13 ad=7.488e-13 ps=1.44e-06 pd=1.13684e-06 sim_w=2.88e-06 m_per_maxw=2.08333 numb_sub_cont=4 nfing=1 $X=76220 $Y=200 $D=21
M31 1 2 1 cpoly_p w=6e-06 l=2e-06 c=8.0712e-14 as=2.1408e-13 ad=7.488e-13 ps=1.44e-06 pd=1.13684e-06 sim_w=2.88e-06 m_per_maxw=2.08333 numb_sub_cont=4 nfing=1 $X=78740 $Y=200 $D=21
M32 1 2 1 cpoly_p w=6e-06 l=2e-06 c=8.0712e-14 as=2.1408e-13 ad=7.488e-13 ps=1.44e-06 pd=1.13684e-06 sim_w=2.88e-06 m_per_maxw=2.08333 numb_sub_cont=4 nfing=1 $X=81260 $Y=200 $D=21
M33 1 2 1 cpoly_p w=6e-06 l=2e-06 c=8.0712e-14 as=2.1408e-13 ad=7.488e-13 ps=1.44e-06 pd=1.13684e-06 sim_w=2.88e-06 m_per_maxw=2.08333 numb_sub_cont=4 nfing=1 $X=83780 $Y=200 $D=21
M34 1 2 1 cpoly_p w=6e-06 l=2e-06 c=8.0712e-14 as=2.1408e-13 ad=7.488e-13 ps=1.44e-06 pd=1.13684e-06 sim_w=2.88e-06 m_per_maxw=2.08333 numb_sub_cont=4 nfing=1 $X=86300 $Y=200 $D=21
M35 1 2 1 cpoly_p w=6e-06 l=2e-06 c=8.0712e-14 as=2.1408e-13 ad=7.488e-13 ps=1.44e-06 pd=1.13684e-06 sim_w=2.88e-06 m_per_maxw=2.08333 numb_sub_cont=4 nfing=1 $X=88820 $Y=200 $D=21
M36 1 2 1 cpoly_p w=6e-06 l=2e-06 c=8.0712e-14 as=2.1408e-13 ad=7.488e-13 ps=1.44e-06 pd=1.13684e-06 sim_w=2.88e-06 m_per_maxw=2.08333 numb_sub_cont=4 nfing=1 $X=91340 $Y=200 $D=21
M37 1 2 1 cpoly_p w=6e-06 l=2e-06 c=8.0712e-14 as=2.1408e-13 ad=7.488e-13 ps=1.44e-06 pd=1.13684e-06 sim_w=2.88e-06 m_per_maxw=2.08333 numb_sub_cont=4 nfing=1 $X=93860 $Y=200 $D=21
M38 1 2 1 cpoly_p w=6e-06 l=2e-06 c=8.0712e-14 as=2.1408e-13 ad=7.488e-13 ps=1.44e-06 pd=1.13684e-06 sim_w=2.88e-06 m_per_maxw=2.08333 numb_sub_cont=4 nfing=1 $X=96380 $Y=200 $D=21
M39 1 2 1 cpoly_p w=6e-06 l=2e-06 c=8.0712e-14 as=2.1408e-13 ad=7.488e-13 ps=1.44e-06 pd=1.13684e-06 sim_w=2.88e-06 m_per_maxw=2.08333 numb_sub_cont=4 nfing=1 $X=98900 $Y=200 $D=21
M40 1 2 1 cpoly_p w=6e-06 l=2e-06 c=8.0712e-14 as=2.1408e-13 ad=7.488e-13 ps=1.44e-06 pd=1.13684e-06 sim_w=2.88e-06 m_per_maxw=2.08333 numb_sub_cont=4 nfing=1 $X=101420 $Y=200 $D=21
M41 1 2 1 cpoly_p w=6e-06 l=2e-06 c=8.0712e-14 as=2.1408e-13 ad=7.488e-13 ps=1.44e-06 pd=1.13684e-06 sim_w=2.88e-06 m_per_maxw=2.08333 numb_sub_cont=4 nfing=1 $X=103940 $Y=200 $D=21
M42 1 2 1 cpoly_p w=6e-06 l=2e-06 c=8.0712e-14 as=2.1408e-13 ad=7.488e-13 ps=1.44e-06 pd=1.13684e-06 sim_w=2.88e-06 m_per_maxw=2.08333 numb_sub_cont=4 nfing=1 $X=106460 $Y=200 $D=21
M43 1 2 1 cpoly_p w=6e-06 l=2e-06 c=8.0712e-14 as=2.1408e-13 ad=7.488e-13 ps=1.44e-06 pd=1.13684e-06 sim_w=2.88e-06 m_per_maxw=2.08333 numb_sub_cont=4 nfing=1 $X=108980 $Y=200 $D=21
M44 1 2 1 cpoly_p w=6e-06 l=2e-06 c=8.0712e-14 as=2.1408e-13 ad=7.488e-13 ps=1.44e-06 pd=1.13684e-06 sim_w=2.88e-06 m_per_maxw=2.08333 numb_sub_cont=4 nfing=1 $X=111500 $Y=200 $D=21
M45 1 2 1 cpoly_p w=6e-06 l=2e-06 c=8.0712e-14 as=2.1408e-13 ad=7.488e-13 ps=1.44e-06 pd=1.13684e-06 sim_w=2.88e-06 m_per_maxw=2.08333 numb_sub_cont=4 nfing=1 $X=114020 $Y=200 $D=21
M46 1 2 1 cpoly_p w=6e-06 l=2e-06 c=8.0712e-14 as=2.1408e-13 ad=7.488e-13 ps=1.44e-06 pd=1.13684e-06 sim_w=2.88e-06 m_per_maxw=2.08333 numb_sub_cont=4 nfing=1 $X=116540 $Y=200 $D=21
M47 1 2 1 cpoly_p w=6e-06 l=2e-06 c=8.0712e-14 as=2.1408e-13 ad=7.488e-13 ps=1.44e-06 pd=1.13684e-06 sim_w=2.88e-06 m_per_maxw=2.08333 numb_sub_cont=4 nfing=1 $X=119060 $Y=200 $D=21
M48 1 2 1 cpoly_p w=6e-06 l=2e-06 c=8.0712e-14 as=2.1408e-13 ad=7.488e-13 ps=1.44e-06 pd=1.13684e-06 sim_w=2.88e-06 m_per_maxw=2.08333 numb_sub_cont=4 nfing=1 $X=121580 $Y=200 $D=21
M49 1 2 1 cpoly_p w=6e-06 l=2e-06 c=8.0712e-14 as=2.1408e-13 ad=7.488e-13 ps=1.44e-06 pd=1.13684e-06 sim_w=2.88e-06 m_per_maxw=2.08333 numb_sub_cont=4 nfing=1 $X=124100 $Y=200 $D=21
M50 1 2 1 cpoly_p w=6e-06 l=2e-06 c=8.0712e-14 as=2.1408e-13 ad=7.488e-13 ps=1.44e-06 pd=1.13684e-06 sim_w=2.88e-06 m_per_maxw=2.08333 numb_sub_cont=4 nfing=1 $X=126620 $Y=200 $D=21
M51 1 2 1 cpoly_p w=6e-06 l=2e-06 c=8.0712e-14 as=2.1408e-13 ad=7.488e-13 ps=1.44e-06 pd=1.13684e-06 sim_w=2.88e-06 m_per_maxw=2.08333 numb_sub_cont=4 nfing=1 $X=129140 $Y=200 $D=21
M52 1 2 1 cpoly_p w=6e-06 l=2e-06 c=8.0712e-14 as=2.1408e-13 ad=7.488e-13 ps=1.44e-06 pd=1.13684e-06 sim_w=2.88e-06 m_per_maxw=2.08333 numb_sub_cont=4 nfing=1 $X=131660 $Y=200 $D=21
M53 1 2 1 cpoly_p w=6e-06 l=2e-06 c=8.0712e-14 as=2.1408e-13 ad=7.488e-13 ps=1.44e-06 pd=1.13684e-06 sim_w=2.88e-06 m_per_maxw=2.08333 numb_sub_cont=4 nfing=1 $X=134180 $Y=200 $D=21
M54 1 2 1 cpoly_p w=6e-06 l=2e-06 c=8.0712e-14 as=2.1408e-13 ad=7.488e-13 ps=1.44e-06 pd=1.13684e-06 sim_w=2.88e-06 m_per_maxw=2.08333 numb_sub_cont=4 nfing=1 $X=136700 $Y=200 $D=21
M55 1 2 1 cpoly_p w=6e-06 l=2e-06 c=8.0712e-14 as=2.1408e-13 ad=7.488e-13 ps=1.44e-06 pd=1.13684e-06 sim_w=2.88e-06 m_per_maxw=2.08333 numb_sub_cont=4 nfing=1 $X=139220 $Y=200 $D=21
M56 1 2 1 cpoly_p w=6e-06 l=2e-06 c=8.0712e-14 as=2.1408e-13 ad=7.488e-13 ps=1.44e-06 pd=1.13684e-06 sim_w=2.88e-06 m_per_maxw=2.08333 numb_sub_cont=4 nfing=1 $X=141740 $Y=200 $D=21
M57 1 2 1 cpoly_p w=6e-06 l=2e-06 c=8.0712e-14 as=2.1408e-13 ad=7.488e-13 ps=1.44e-06 pd=1.13684e-06 sim_w=2.88e-06 m_per_maxw=2.08333 numb_sub_cont=4 nfing=1 $X=144260 $Y=200 $D=21
M58 1 2 1 cpoly_p w=6e-06 l=2e-06 c=8.0712e-14 as=2.1408e-13 ad=7.488e-13 ps=1.44e-06 pd=1.13684e-06 sim_w=2.88e-06 m_per_maxw=2.08333 numb_sub_cont=4 nfing=1 $X=146780 $Y=200 $D=21
M59 1 2 1 cpoly_p w=6e-06 l=2e-06 c=8.0712e-14 as=2.1408e-13 ad=7.488e-13 ps=1.44e-06 pd=1.13684e-06 sim_w=2.88e-06 m_per_maxw=2.08333 numb_sub_cont=4 nfing=1 $X=149300 $Y=200 $D=21
M60 1 2 1 cpoly_p w=6e-06 l=2e-06 c=8.0712e-14 as=2.1408e-13 ad=7.488e-13 ps=1.44e-06 pd=1.13684e-06 sim_w=2.88e-06 m_per_maxw=2.08333 numb_sub_cont=4 nfing=1 $X=151820 $Y=200 $D=21
M61 1 2 1 cpoly_p w=6e-06 l=2e-06 c=8.0712e-14 as=2.1408e-13 ad=7.488e-13 ps=1.44e-06 pd=1.13684e-06 sim_w=2.88e-06 m_per_maxw=2.08333 numb_sub_cont=4 nfing=1 $X=154340 $Y=200 $D=21
M62 1 2 1 cpoly_p w=6e-06 l=2e-06 c=8.0712e-14 as=2.1408e-13 ad=7.488e-13 ps=1.44e-06 pd=1.13684e-06 sim_w=2.88e-06 m_per_maxw=2.08333 numb_sub_cont=4 nfing=1 $X=156860 $Y=200 $D=21
M63 1 2 1 cpoly_p w=6e-06 l=2e-06 c=8.0712e-14 as=2.1408e-13 ad=7.488e-13 ps=1.44e-06 pd=1.13684e-06 sim_w=2.88e-06 m_per_maxw=2.08333 numb_sub_cont=4 nfing=1 $X=159380 $Y=200 $D=21
M64 1 2 1 cpoly_p w=6e-06 l=2e-06 c=8.0712e-14 as=2.1408e-13 ad=7.488e-13 ps=1.44e-06 pd=1.13684e-06 sim_w=2.88e-06 m_per_maxw=2.08333 numb_sub_cont=4 nfing=1 $X=161900 $Y=200 $D=21
M65 1 2 1 cpoly_p w=6e-06 l=2e-06 c=8.0712e-14 as=2.1408e-13 ad=7.488e-13 ps=1.44e-06 pd=1.13684e-06 sim_w=2.88e-06 m_per_maxw=2.08333 numb_sub_cont=4 nfing=1 $X=164420 $Y=200 $D=21
M66 1 2 1 cpoly_p w=6e-06 l=2e-06 c=8.0712e-14 as=2.1408e-13 ad=7.488e-13 ps=1.44e-06 pd=1.13684e-06 sim_w=2.88e-06 m_per_maxw=2.08333 numb_sub_cont=4 nfing=1 $X=166940 $Y=200 $D=21
M67 1 2 1 cpoly_p w=6e-06 l=2e-06 c=8.0712e-14 as=2.1408e-13 ad=7.488e-13 ps=1.44e-06 pd=1.13684e-06 sim_w=2.88e-06 m_per_maxw=2.08333 numb_sub_cont=4 nfing=1 $X=169460 $Y=200 $D=21
M68 1 2 1 cpoly_p w=6e-06 l=2e-06 c=8.0712e-14 as=2.1408e-13 ad=7.488e-13 ps=1.44e-06 pd=1.13684e-06 sim_w=2.88e-06 m_per_maxw=2.08333 numb_sub_cont=4 nfing=1 $X=171980 $Y=200 $D=21
M69 1 2 1 cpoly_p w=6e-06 l=2e-06 c=8.0712e-14 as=2.1408e-13 ad=7.488e-13 ps=1.44e-06 pd=1.13684e-06 sim_w=2.88e-06 m_per_maxw=2.08333 numb_sub_cont=4 nfing=1 $X=174500 $Y=200 $D=21
M70 1 2 1 cpoly_p w=6e-06 l=2e-06 c=8.0712e-14 as=2.1408e-13 ad=7.488e-13 ps=1.44e-06 pd=1.13684e-06 sim_w=2.88e-06 m_per_maxw=2.08333 numb_sub_cont=4 nfing=1 $X=177020 $Y=200 $D=21
M71 1 2 1 cpoly_p w=6e-06 l=2e-06 c=8.0712e-14 as=2.1408e-13 ad=7.488e-13 ps=1.44e-06 pd=1.13684e-06 sim_w=2.88e-06 m_per_maxw=2.08333 numb_sub_cont=4 nfing=1 $X=179540 $Y=200 $D=21
M72 1 2 1 cpoly_p w=6e-06 l=2e-06 c=8.0712e-14 as=2.1408e-13 ad=7.488e-13 ps=1.44e-06 pd=1.13684e-06 sim_w=2.88e-06 m_per_maxw=2.08333 numb_sub_cont=4 nfing=1 $X=182060 $Y=200 $D=21
M73 1 2 1 cpoly_p w=6e-06 l=2e-06 c=8.0712e-14 as=2.1408e-13 ad=7.488e-13 ps=1.44e-06 pd=1.13684e-06 sim_w=2.88e-06 m_per_maxw=2.08333 numb_sub_cont=4 nfing=1 $X=184580 $Y=200 $D=21
M74 1 2 1 cpoly_p w=6e-06 l=2e-06 c=8.0712e-14 as=2.1408e-13 ad=7.488e-13 ps=1.44e-06 pd=1.13684e-06 sim_w=2.88e-06 m_per_maxw=2.08333 numb_sub_cont=4 nfing=1 $X=187100 $Y=200 $D=21
M75 1 2 1 cpoly_p w=6e-06 l=2e-06 c=8.0712e-14 as=2.1408e-13 ad=7.488e-13 ps=1.44e-06 pd=1.13684e-06 sim_w=2.88e-06 m_per_maxw=2.08333 numb_sub_cont=4 nfing=1 $X=189620 $Y=200 $D=21
M76 1 2 1 cpoly_p w=6e-06 l=2e-06 c=8.0712e-14 as=2.1408e-13 ad=7.488e-13 ps=1.44e-06 pd=1.13684e-06 sim_w=2.88e-06 m_per_maxw=2.08333 numb_sub_cont=4 nfing=1 $X=192140 $Y=200 $D=21
M77 1 2 1 cpoly_p w=6e-06 l=2e-06 c=8.0712e-14 as=2.1408e-13 ad=7.488e-13 ps=1.44e-06 pd=1.13684e-06 sim_w=2.88e-06 m_per_maxw=2.08333 numb_sub_cont=4 nfing=1 $X=194660 $Y=200 $D=21
M78 1 2 1 cpoly_p w=6e-06 l=2e-06 c=8.0712e-14 as=2.1408e-13 ad=7.488e-13 ps=1.44e-06 pd=1.13684e-06 sim_w=2.88e-06 m_per_maxw=2.08333 numb_sub_cont=4 nfing=1 $X=197180 $Y=200 $D=21
M79 1 2 1 cpoly_p w=6e-06 l=2e-06 c=8.0712e-14 as=1.68e-13 ad=7.488e-13 ps=1.44e-06 pd=1.13684e-06 sim_w=2.88e-06 m_per_maxw=2.08333 numb_sub_cont=4 nfing=1 $X=199700 $Y=200 $D=21
.ENDS
***************************************
.SUBCKT rppoly_CDNS_5887047866532 1 2
** N=2 EP=2 IP=0 FDC=1
R0 1 2 18955.3 L=0.00020234 W=3.44e-06 m=1 $[rppoly] $X=0 $Y=0 $D=19
.ENDS
***************************************
.SUBCKT cpoly_p_CDNS_5887047866534 1 2
** N=2 EP=2 IP=0 FDC=4
M0 1 2 1 cpoly_p w=1e-05 l=2e-06 c=1.28502e-13 as=1.3536e-13 ad=7.488e-13 ps=1.44e-06 pd=1.19008e-06 sim_w=2.88e-06 m_per_maxw=3.47222 numb_sub_cont=5 nfing=1 $X=620 $Y=200 $D=21
M1 1 2 1 cpoly_p w=1e-05 l=2e-06 c=1.28502e-13 as=1.71648e-13 ad=7.488e-13 ps=1.44e-06 pd=1.19008e-06 sim_w=2.88e-06 m_per_maxw=3.47222 numb_sub_cont=5 nfing=1 $X=3140 $Y=200 $D=21
M2 1 2 1 cpoly_p w=1e-05 l=2e-06 c=1.28502e-13 as=1.71648e-13 ad=7.488e-13 ps=1.44e-06 pd=1.19008e-06 sim_w=2.88e-06 m_per_maxw=3.47222 numb_sub_cont=5 nfing=1 $X=5660 $Y=200 $D=21
M3 1 2 1 cpoly_p w=1e-05 l=2e-06 c=1.28502e-13 as=1.3536e-13 ad=7.488e-13 ps=1.44e-06 pd=1.19008e-06 sim_w=2.88e-06 m_per_maxw=3.47222 numb_sub_cont=5 nfing=1 $X=8180 $Y=200 $D=21
.ENDS
***************************************
.SUBCKT ICV_34 1 2
** N=2 EP=2 IP=4 FDC=8
X0 1 2 cpoly_p_CDNS_5887047866534 $T=0 0 0 0 $X=0 $Y=0
X1 1 2 cpoly_p_CDNS_5887047866534 $T=10760 0 0 0 $X=10760 $Y=0
.ENDS
***************************************
.SUBCKT PAD_Clamp_160 gnd! vdd!
** N=6 EP=2 IP=372 FDC=1405
M0 5 4 vdd! vdd! pmos_a L=2.4e-07 W=4e-06 AD=1.84e-12 AS=1.4e-13 PD=4.6e-06 PS=2.3e-06 w_cont=6e-07 nfing=1 mmm=1 $X=34040 $Y=45280 $D=5
M1 5 4 vdd! vdd! pmos_a L=2.4e-07 W=4e-06 AD=1.84e-12 AS=1.4e-13 PD=4.6e-06 PS=2.3e-06 w_cont=6e-07 nfing=1 mmm=1 $X=34040 $Y=155280 $D=5
M2 5 4 vdd! vdd! pmos_a L=2.4e-07 W=4e-06 AD=1.84e-12 AS=1.4e-13 PD=4.6e-06 PS=2.3e-06 w_cont=6e-07 nfing=1 mmm=1 $X=39540 $Y=45280 $D=5
M3 5 4 vdd! vdd! pmos_a L=2.4e-07 W=4e-06 AD=1.84e-12 AS=1.4e-13 PD=4.6e-06 PS=2.3e-06 w_cont=6e-07 nfing=1 mmm=1 $X=39540 $Y=155280 $D=5
M4 5 4 vdd! vdd! pmos_a L=2.4e-07 W=4e-06 AD=1.84e-12 AS=1.4e-13 PD=4.6e-06 PS=2.3e-06 w_cont=6e-07 nfing=1 mmm=1 $X=53540 $Y=45280 $D=5
M5 5 4 vdd! vdd! pmos_a L=2.4e-07 W=4e-06 AD=1.84e-12 AS=1.4e-13 PD=4.6e-06 PS=2.3e-06 w_cont=6e-07 nfing=1 mmm=1 $X=53540 $Y=155280 $D=5
M6 5 4 vdd! vdd! pmos_a L=2.4e-07 W=4e-06 AD=1.84e-12 AS=1.4e-13 PD=4.6e-06 PS=2.3e-06 w_cont=6e-07 nfing=1 mmm=1 $X=62040 $Y=45280 $D=5
M7 5 4 vdd! vdd! pmos_a L=2.4e-07 W=4e-06 AD=1.84e-12 AS=1.4e-13 PD=4.6e-06 PS=2.3e-06 w_cont=6e-07 nfing=1 mmm=1 $X=62040 $Y=155280 $D=5
M8 4 3 vdd! vdd! pmos_a L=2.4e-07 W=4e-06 AD=1.84e-12 AS=1.4e-13 PD=4.6e-06 PS=2.3e-06 w_cont=6e-07 nfing=1 mmm=1 $X=68740 $Y=105760 $D=5
M9 4 3 vdd! vdd! pmos_a L=2.4e-07 W=4e-06 AD=1.84e-12 AS=1.4e-13 PD=4.6e-06 PS=2.3e-06 w_cont=6e-07 nfing=1 mmm=1 $X=68740 $Y=115000 $D=5
M10 4 3 vdd! vdd! pmos_a L=2.4e-07 W=4e-06 AD=1.84e-12 AS=1.4e-13 PD=4.6e-06 PS=2.3e-06 w_cont=6e-07 nfing=1 mmm=1 $X=68740 $Y=124400 $D=5
M11 4 3 vdd! vdd! pmos_a L=2.4e-07 W=4e-06 AD=1.84e-12 AS=1.4e-13 PD=4.6e-06 PS=2.3e-06 w_cont=6e-07 nfing=1 mmm=1 $X=68740 $Y=133920 $D=5
M12 4 3 vdd! vdd! pmos_a L=2.4e-07 W=4e-06 AD=1.84e-12 AS=1.4e-13 PD=4.6e-06 PS=2.3e-06 w_cont=6e-07 nfing=1 mmm=1 $X=81880 $Y=105760 $D=5
M13 4 3 vdd! vdd! pmos_a L=2.4e-07 W=4e-06 AD=1.84e-12 AS=1.4e-13 PD=4.6e-06 PS=2.3e-06 w_cont=6e-07 nfing=1 mmm=1 $X=81880 $Y=115000 $D=5
M14 4 3 vdd! vdd! pmos_a L=2.4e-07 W=4e-06 AD=1.84e-12 AS=1.4e-13 PD=4.6e-06 PS=2.3e-06 w_cont=6e-07 nfing=1 mmm=1 $X=81880 $Y=124400 $D=5
M15 4 3 vdd! vdd! pmos_a L=2.4e-07 W=4e-06 AD=1.84e-12 AS=1.4e-13 PD=4.6e-06 PS=2.3e-06 w_cont=6e-07 nfing=1 mmm=1 $X=81880 $Y=133920 $D=5
M16 5 4 vdd! vdd! pmos_a L=2.4e-07 W=4e-06 AD=1.84e-12 AS=1.4e-13 PD=4.6e-06 PS=2.3e-06 w_cont=6e-07 nfing=1 mmm=1 $X=90040 $Y=45280 $D=5
M17 5 4 vdd! vdd! pmos_a L=2.4e-07 W=4e-06 AD=1.84e-12 AS=1.4e-13 PD=4.6e-06 PS=2.3e-06 w_cont=6e-07 nfing=1 mmm=1 $X=90040 $Y=155280 $D=5
M18 5 4 vdd! vdd! pmos_a L=2.4e-07 W=4e-06 AD=1.84e-12 AS=1.4e-13 PD=4.6e-06 PS=2.3e-06 w_cont=6e-07 nfing=1 mmm=1 $X=95540 $Y=45280 $D=5
M19 5 4 vdd! vdd! pmos_a L=2.4e-07 W=4e-06 AD=1.84e-12 AS=1.4e-13 PD=4.6e-06 PS=2.3e-06 w_cont=6e-07 nfing=1 mmm=1 $X=95540 $Y=155280 $D=5
M20 5 4 vdd! vdd! pmos_a L=2.4e-07 W=4e-06 AD=1.84e-12 AS=1.4e-13 PD=4.6e-06 PS=2.3e-06 w_cont=6e-07 nfing=1 mmm=1 $X=109540 $Y=45280 $D=5
M21 5 4 vdd! vdd! pmos_a L=2.4e-07 W=4e-06 AD=1.84e-12 AS=1.4e-13 PD=4.6e-06 PS=2.3e-06 w_cont=6e-07 nfing=1 mmm=1 $X=109540 $Y=155280 $D=5
M22 5 4 vdd! vdd! pmos_a L=2.4e-07 W=4e-06 AD=1.84e-12 AS=1.4e-13 PD=4.6e-06 PS=2.3e-06 w_cont=6e-07 nfing=1 mmm=1 $X=118040 $Y=45280 $D=5
M23 5 4 vdd! vdd! pmos_a L=2.4e-07 W=4e-06 AD=1.84e-12 AS=1.4e-13 PD=4.6e-06 PS=2.3e-06 w_cont=6e-07 nfing=1 mmm=1 $X=118040 $Y=155280 $D=5
X24 gnd! vdd! cpoly_p_CDNS_58870478665105 $T=1240 420500 0 0 $X=1240 $Y=420500
X25 vdd! gnd! cpoly_n_CDNS_58870478665104 $T=1220 433340 0 0 $X=1220 $Y=433340
X26 gnd! vdd! cpoly_p_CDNS_5887047866536 $T=17580 220 0 90 $X=9580 $Y=220
X27 gnd! vdd! cpoly_p_CDNS_5887047866536 $T=130740 220 0 90 $X=122740 $Y=220
X28 vdd! gnd! cpoly_n_CDNS_5887047866529 $T=26760 0 0 90 $X=19260 $Y=0
X29 vdd! gnd! cpoly_n_CDNS_5887047866529 $T=144860 0 0 90 $X=137360 $Y=0
X54 gnd! vdd! 5 nmos_io_a_CDNS_5887047866531 $T=31960 260 0 0 $X=31960 $Y=160
X55 gnd! vdd! 5 nmos_io_a_CDNS_5887047866531 $T=31960 25720 0 0 $X=31960 $Y=25620
X56 gnd! vdd! 5 nmos_io_a_CDNS_5887047866531 $T=31960 55060 0 0 $X=31960 $Y=54960
X57 gnd! vdd! 5 nmos_io_a_CDNS_5887047866531 $T=31960 82460 0 0 $X=31960 $Y=82360
X58 gnd! vdd! 5 nmos_io_a_CDNS_5887047866531 $T=31960 109860 0 0 $X=31960 $Y=109760
X59 gnd! vdd! 5 nmos_io_a_CDNS_5887047866531 $T=31960 137260 0 0 $X=31960 $Y=137160
X60 gnd! vdd! 5 nmos_io_a_CDNS_5887047866531 $T=31960 164660 0 0 $X=31960 $Y=164560
X61 gnd! vdd! 5 nmos_io_a_CDNS_5887047866531 $T=31960 190400 0 0 $X=31960 $Y=190300
X62 gnd! vdd! 5 nmos_io_a_CDNS_5887047866531 $T=41860 260 1 180 $X=38960 $Y=160
X63 gnd! vdd! 5 nmos_io_a_CDNS_5887047866531 $T=41860 25720 1 180 $X=38960 $Y=25620
X64 gnd! vdd! 5 nmos_io_a_CDNS_5887047866531 $T=41860 55060 1 180 $X=38960 $Y=54960
X65 gnd! vdd! 5 nmos_io_a_CDNS_5887047866531 $T=41860 82460 1 180 $X=38960 $Y=82360
X66 gnd! vdd! 5 nmos_io_a_CDNS_5887047866531 $T=41860 109860 1 180 $X=38960 $Y=109760
X67 gnd! vdd! 5 nmos_io_a_CDNS_5887047866531 $T=41860 137260 1 180 $X=38960 $Y=137160
X68 gnd! vdd! 5 nmos_io_a_CDNS_5887047866531 $T=41860 164660 1 180 $X=38960 $Y=164560
X69 gnd! vdd! 5 nmos_io_a_CDNS_5887047866531 $T=41860 190400 1 180 $X=38960 $Y=190300
X70 gnd! vdd! 5 nmos_io_a_CDNS_5887047866531 $T=45960 260 0 0 $X=45960 $Y=160
X71 gnd! vdd! 5 nmos_io_a_CDNS_5887047866531 $T=45960 25720 0 0 $X=45960 $Y=25620
X72 gnd! vdd! 5 nmos_io_a_CDNS_5887047866531 $T=45960 55060 0 0 $X=45960 $Y=54960
X73 gnd! vdd! 5 nmos_io_a_CDNS_5887047866531 $T=45960 82460 0 0 $X=45960 $Y=82360
X74 gnd! vdd! 5 nmos_io_a_CDNS_5887047866531 $T=45960 109860 0 0 $X=45960 $Y=109760
X75 gnd! vdd! 5 nmos_io_a_CDNS_5887047866531 $T=45960 137260 0 0 $X=45960 $Y=137160
X76 gnd! vdd! 5 nmos_io_a_CDNS_5887047866531 $T=45960 164660 0 0 $X=45960 $Y=164560
X77 gnd! vdd! 5 nmos_io_a_CDNS_5887047866531 $T=45960 190400 0 0 $X=45960 $Y=190300
X78 gnd! vdd! 5 nmos_io_a_CDNS_5887047866531 $T=55860 260 1 180 $X=52960 $Y=160
X79 gnd! vdd! 5 nmos_io_a_CDNS_5887047866531 $T=55860 25720 1 180 $X=52960 $Y=25620
X80 gnd! vdd! 5 nmos_io_a_CDNS_5887047866531 $T=55860 55060 1 180 $X=52960 $Y=54960
X81 gnd! vdd! 5 nmos_io_a_CDNS_5887047866531 $T=55860 82460 1 180 $X=52960 $Y=82360
X82 gnd! vdd! 5 nmos_io_a_CDNS_5887047866531 $T=55860 109860 1 180 $X=52960 $Y=109760
X83 gnd! vdd! 5 nmos_io_a_CDNS_5887047866531 $T=55860 137260 1 180 $X=52960 $Y=137160
X84 gnd! vdd! 5 nmos_io_a_CDNS_5887047866531 $T=55860 164660 1 180 $X=52960 $Y=164560
X85 gnd! vdd! 5 nmos_io_a_CDNS_5887047866531 $T=55860 190400 1 180 $X=52960 $Y=190300
X86 gnd! vdd! 5 nmos_io_a_CDNS_5887047866531 $T=59960 260 0 0 $X=59960 $Y=160
X87 gnd! vdd! 5 nmos_io_a_CDNS_5887047866531 $T=59960 25720 0 0 $X=59960 $Y=25620
X88 gnd! vdd! 5 nmos_io_a_CDNS_5887047866531 $T=59960 55060 0 0 $X=59960 $Y=54960
X89 gnd! vdd! 5 nmos_io_a_CDNS_5887047866531 $T=59960 82460 0 0 $X=59960 $Y=82360
X90 gnd! vdd! 5 nmos_io_a_CDNS_5887047866531 $T=59960 109860 0 0 $X=59960 $Y=109760
X91 gnd! vdd! 5 nmos_io_a_CDNS_5887047866531 $T=59960 137260 0 0 $X=59960 $Y=137160
X92 gnd! vdd! 5 nmos_io_a_CDNS_5887047866531 $T=59960 164660 0 0 $X=59960 $Y=164560
X93 gnd! vdd! 5 nmos_io_a_CDNS_5887047866531 $T=59960 190400 0 0 $X=59960 $Y=190300
X94 gnd! vdd! 5 nmos_io_a_CDNS_5887047866531 $T=87960 260 0 0 $X=87960 $Y=160
X95 gnd! vdd! 5 nmos_io_a_CDNS_5887047866531 $T=87960 25660 0 0 $X=87960 $Y=25560
X96 gnd! vdd! 5 nmos_io_a_CDNS_5887047866531 $T=87960 55060 0 0 $X=87960 $Y=54960
X97 gnd! vdd! 5 nmos_io_a_CDNS_5887047866531 $T=87960 82460 0 0 $X=87960 $Y=82360
X98 gnd! vdd! 5 nmos_io_a_CDNS_5887047866531 $T=87960 109860 0 0 $X=87960 $Y=109760
X99 gnd! vdd! 5 nmos_io_a_CDNS_5887047866531 $T=87960 137260 0 0 $X=87960 $Y=137160
X100 gnd! vdd! 5 nmos_io_a_CDNS_5887047866531 $T=87960 164660 0 0 $X=87960 $Y=164560
X101 gnd! vdd! 5 nmos_io_a_CDNS_5887047866531 $T=87960 190400 0 0 $X=87960 $Y=190300
X102 gnd! vdd! 5 nmos_io_a_CDNS_5887047866531 $T=97860 260 1 180 $X=94960 $Y=160
X103 gnd! vdd! 5 nmos_io_a_CDNS_5887047866531 $T=97860 25660 1 180 $X=94960 $Y=25560
X104 gnd! vdd! 5 nmos_io_a_CDNS_5887047866531 $T=97860 55060 1 180 $X=94960 $Y=54960
X105 gnd! vdd! 5 nmos_io_a_CDNS_5887047866531 $T=97860 82460 1 180 $X=94960 $Y=82360
X106 gnd! vdd! 5 nmos_io_a_CDNS_5887047866531 $T=97860 109860 1 180 $X=94960 $Y=109760
X107 gnd! vdd! 5 nmos_io_a_CDNS_5887047866531 $T=97860 137260 1 180 $X=94960 $Y=137160
X108 gnd! vdd! 5 nmos_io_a_CDNS_5887047866531 $T=97860 164660 1 180 $X=94960 $Y=164560
X109 gnd! vdd! 5 nmos_io_a_CDNS_5887047866531 $T=97860 190400 1 180 $X=94960 $Y=190300
X110 gnd! vdd! 5 nmos_io_a_CDNS_5887047866531 $T=101960 260 0 0 $X=101960 $Y=160
X111 gnd! vdd! 5 nmos_io_a_CDNS_5887047866531 $T=101960 25660 0 0 $X=101960 $Y=25560
X112 gnd! vdd! 5 nmos_io_a_CDNS_5887047866531 $T=101960 55060 0 0 $X=101960 $Y=54960
X113 gnd! vdd! 5 nmos_io_a_CDNS_5887047866531 $T=101960 82460 0 0 $X=101960 $Y=82360
X114 gnd! vdd! 5 nmos_io_a_CDNS_5887047866531 $T=101960 109860 0 0 $X=101960 $Y=109760
X115 gnd! vdd! 5 nmos_io_a_CDNS_5887047866531 $T=101960 137260 0 0 $X=101960 $Y=137160
X116 gnd! vdd! 5 nmos_io_a_CDNS_5887047866531 $T=101960 164660 0 0 $X=101960 $Y=164560
X117 gnd! vdd! 5 nmos_io_a_CDNS_5887047866531 $T=101960 190400 0 0 $X=101960 $Y=190300
X118 gnd! vdd! 5 nmos_io_a_CDNS_5887047866531 $T=111860 260 1 180 $X=108960 $Y=160
X119 gnd! vdd! 5 nmos_io_a_CDNS_5887047866531 $T=111860 25660 1 180 $X=108960 $Y=25560
X120 gnd! vdd! 5 nmos_io_a_CDNS_5887047866531 $T=111860 55060 1 180 $X=108960 $Y=54960
X121 gnd! vdd! 5 nmos_io_a_CDNS_5887047866531 $T=111860 82460 1 180 $X=108960 $Y=82360
X122 gnd! vdd! 5 nmos_io_a_CDNS_5887047866531 $T=111860 109860 1 180 $X=108960 $Y=109760
X123 gnd! vdd! 5 nmos_io_a_CDNS_5887047866531 $T=111860 137260 1 180 $X=108960 $Y=137160
X124 gnd! vdd! 5 nmos_io_a_CDNS_5887047866531 $T=111860 164660 1 180 $X=108960 $Y=164560
X125 gnd! vdd! 5 nmos_io_a_CDNS_5887047866531 $T=111860 190400 1 180 $X=108960 $Y=190300
X126 gnd! vdd! 5 nmos_io_a_CDNS_5887047866531 $T=115960 260 0 0 $X=115960 $Y=160
X127 gnd! vdd! 5 nmos_io_a_CDNS_5887047866531 $T=115960 25660 0 0 $X=115960 $Y=25560
X128 gnd! vdd! 5 nmos_io_a_CDNS_5887047866531 $T=115960 55060 0 0 $X=115960 $Y=54960
X129 gnd! vdd! 5 nmos_io_a_CDNS_5887047866531 $T=115960 82460 0 0 $X=115960 $Y=82360
X130 gnd! vdd! 5 nmos_io_a_CDNS_5887047866531 $T=115960 109860 0 0 $X=115960 $Y=109760
X131 gnd! vdd! 5 nmos_io_a_CDNS_5887047866531 $T=115960 137260 0 0 $X=115960 $Y=137160
X132 gnd! vdd! 5 nmos_io_a_CDNS_5887047866531 $T=115960 164660 0 0 $X=115960 $Y=164560
X133 gnd! vdd! 5 nmos_io_a_CDNS_5887047866531 $T=115960 190400 0 0 $X=115960 $Y=190300
X134 vdd! gnd! cpoly_n_CDNS_5887047866535 $T=56340 211680 0 90 $X=48840 $Y=211680
X135 vdd! gnd! cpoly_n_CDNS_5887047866535 $T=85800 211680 0 90 $X=78300 $Y=211680
X136 vdd! gnd! cpoly_n_CDNS_5887047866535 $T=115260 211680 0 90 $X=107760 $Y=211680
X137 gnd! 5 4 nmos_a_CDNS_5887047866530 $T=45960 43580 0 0 $X=45960 $Y=43580
X138 gnd! 5 4 nmos_a_CDNS_5887047866530 $T=45960 155080 0 0 $X=45960 $Y=155080
X139 gnd! 4 3 nmos_a_CDNS_5887047866530 $T=69600 86980 1 180 $X=68160 $Y=86980
X140 gnd! 4 3 nmos_a_CDNS_5887047866530 $T=69600 94920 1 180 $X=68160 $Y=94920
X141 gnd! 4 3 nmos_a_CDNS_5887047866530 $T=81260 86980 0 0 $X=81260 $Y=86980
X142 gnd! 4 3 nmos_a_CDNS_5887047866530 $T=81260 94940 0 0 $X=81260 $Y=94940
X143 gnd! 5 4 nmos_a_CDNS_5887047866530 $T=101960 43580 0 0 $X=101960 $Y=43580
X144 gnd! 5 4 nmos_a_CDNS_5887047866530 $T=101960 155080 0 0 $X=101960 $Y=155080
X145 gnd! vdd! cpoly_p_CDNS_5887047866528 $T=42220 211900 0 90 $X=34220 $Y=211900
X146 gnd! vdd! cpoly_p_CDNS_5887047866528 $T=71680 211900 0 90 $X=63680 $Y=211900
X147 gnd! vdd! cpoly_p_CDNS_5887047866528 $T=101140 211900 0 90 $X=93140 $Y=211900
X148 gnd! 3 rppoly_CDNS_5887047866532 $T=86920 204240 1 270 $X=83180 $Y=1140
X149 3 vdd! cpoly_p_CDNS_5887047866534 $T=69020 140 1 90 $X=69020 $Y=140
X150 3 vdd! cpoly_p_CDNS_5887047866534 $T=69020 75480 1 90 $X=69020 $Y=75480
X151 3 vdd! ICV_34 $T=69020 10920 1 90 $X=69020 $Y=10920
X152 3 vdd! ICV_34 $T=69020 32440 1 90 $X=69020 $Y=32440
X153 3 vdd! ICV_34 $T=69020 53960 1 90 $X=69020 $Y=53960
.ENDS
***************************************
.SUBCKT ICV_35
** N=2 EP=0 IP=4 FDC=0
.ENDS
***************************************
.SUBCKT ICV_36 1 2
** N=2 EP=2 IP=4 FDC=4
D0 2 1 dn PJ=0.00041 m=1 $X=2720 $Y=0 $D=8
D1 2 1 dn PJ=0.00041 m=1 $X=7720 $Y=0 $D=8
D2 2 1 dn PJ=0.00041 m=1 $X=-460 $Y=0 $D=9
D3 2 1 dn PJ=0.00041 m=1 $X=4540 $Y=0 $D=9
.ENDS
***************************************
.SUBCKT ICV_37 1 2
** N=2 EP=2 IP=4 FDC=8
X0 1 2 ICV_36 $T=0 0 0 0 $X=-640 $Y=-300
X1 1 2 ICV_36 $T=10000 0 0 0 $X=9360 $Y=-300
.ENDS
***************************************
.SUBCKT VDD_Core vdd! gnd!
** N=6 EP=2 IP=16 FDC=115
D0 gnd! vdd! dn PJ=0.00041 m=1 $X=94280 $Y=-99700 $D=9
X1 vdd! gnd! cpoly_n_CDNS_588704786651 $T=520 333340 0 0 $X=520 $Y=333340
X2 gnd! vdd! cpoly_p_CDNS_588704786650 $T=520 320500 0 0 $X=520 $Y=320500
X4 vdd! gnd! ICV_36 $T=84740 -99700 0 0 $X=84100 $Y=-100000
X5 vdd! gnd! ICV_37 $T=4740 -99700 0 0 $X=4100 $Y=-100000
X6 vdd! gnd! ICV_37 $T=24740 -99700 0 0 $X=24100 $Y=-100000
X7 vdd! gnd! ICV_37 $T=44740 -99700 0 0 $X=44100 $Y=-100000
X8 vdd! gnd! ICV_37 $T=64740 -99700 0 0 $X=64100 $Y=-100000
.ENDS
***************************************
.SUBCKT ICV_38 1 2 3 4 6 7 8 9 10 11 12 13 14
** N=14 EP=13 IP=20 FDC=5490
X0 1 2 3 4 7 6 10 9 13 ICV_30 $T=-300000 0 0 0 $X=-405000 $Y=-136000
X1 1 2 3 4 7 8 12 11 14 ICV_30 $T=0 0 0 0 $X=-105000 $Y=-136000
.ENDS
***************************************
.SUBCKT ICV_39 1 2
** N=5 EP=2 IP=8 FDC=3576
X0 1 2 Fill_Block_8Kx8 $T=0 0 0 0 $X=-360 $Y=-320
X1 1 2 Fill_Block_8Kx8 $T=440480 0 0 0 $X=440120 $Y=-320
.ENDS
***************************************
.SUBCKT ICV_40 1 2
** N=2 EP=2 IP=2 FDC=78
X0 1 2 cpoly_n_CDNS_5887047866527 $T=0 0 0 0 $X=0 $Y=0
.ENDS
***************************************
.SUBCKT ICV_41 1 2
** N=2 EP=2 IP=2 FDC=78
X0 1 2 cpoly_p_CDNS_5887047866533 $T=0 0 0 0 $X=0 $Y=0
.ENDS
***************************************
.SUBCKT ICV_42 1 2
** N=2 EP=2 IP=2 FDC=80
X0 1 2 cpoly_p_CDNS_5887047866528 $T=0 0 0 0 $X=0 $Y=0
.ENDS
***************************************
.SUBCKT ICV_43 1 2
** N=2 EP=2 IP=2 FDC=164
X0 1 2 cpoly_p_CDNS_5887047866536 $T=0 0 0 0 $X=0 $Y=0
.ENDS
***************************************
.SUBCKT ICV_44 1 2
** N=2 EP=2 IP=2 FDC=164
X0 1 2 cpoly_p_CDNS_5887047866536 $T=0 0 0 0 $X=0 $Y=0
.ENDS
***************************************
.SUBCKT ICV_45 1 2
** N=2 EP=2 IP=2 FDC=164
X0 1 2 cpoly_p_CDNS_5887047866536 $T=0 0 0 0 $X=0 $Y=0
.ENDS
***************************************
.SUBCKT ICV_46 1 2
** N=2 EP=2 IP=2 FDC=164
X0 1 2 cpoly_p_CDNS_5887047866536 $T=0 0 0 0 $X=0 $Y=0
.ENDS
***************************************
.SUBCKT ICV_47 1 2
** N=2 EP=2 IP=2 FDC=164
X0 1 2 cpoly_p_CDNS_5887047866536 $T=0 0 0 0 $X=0 $Y=0
.ENDS
***************************************
.SUBCKT ICV_48 1 2
** N=2 EP=2 IP=2 FDC=164
X0 2 1 cpoly_n_CDNS_5887047866529 $T=0 0 0 0 $X=0 $Y=0
.ENDS
***************************************
.SUBCKT ICV_49 1 2
** N=2 EP=2 IP=2 FDC=164
X0 2 1 cpoly_n_CDNS_5887047866529 $T=0 0 0 0 $X=0 $Y=0
.ENDS
***************************************
.SUBCKT ICV_50 1 2
** N=2 EP=2 IP=2 FDC=164
X0 2 1 cpoly_n_CDNS_5887047866529 $T=0 0 0 0 $X=0 $Y=0
.ENDS
***************************************
.SUBCKT ICV_51 1 2
** N=2 EP=2 IP=2 FDC=164
X0 2 1 cpoly_n_CDNS_5887047866529 $T=0 0 0 0 $X=0 $Y=0
.ENDS
***************************************
.SUBCKT ICV_52 1 2
** N=2 EP=2 IP=2 FDC=164
X0 2 1 cpoly_n_CDNS_5887047866529 $T=0 0 0 0 $X=0 $Y=0
.ENDS
***************************************
.SUBCKT ICV_53
** N=4 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT ICV_54
** N=2 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT ICV_55
** N=2 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT ICV_56
** N=2 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT ICV_57
** N=3 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT ICV_58 1 2 5
** N=5 EP=3 IP=14 FDC=84
X0 2 1 5 nmos_io_a_CDNS_5887047866531 $T=190400 -165660 0 270 $X=190300 $Y=-168560
X1 2 1 5 nmos_io_a_CDNS_5887047866531 $T=190400 -161560 1 90 $X=190300 $Y=-161560
X2 2 1 5 nmos_io_a_CDNS_5887047866531 $T=190400 -151660 0 270 $X=190300 $Y=-154560
X3 2 1 5 nmos_io_a_CDNS_5887047866531 $T=190400 -147560 1 90 $X=190300 $Y=-147560
X4 1 2 cpoly_n_CDNS_5887047866535 $T=211680 -164960 0 0 $X=211680 $Y=-164960
.ENDS
***************************************
.SUBCKT ICV_59 1 2 3 4
** N=4 EP=4 IP=36 FDC=12
M0 3 2 1 1 pmos_a L=2.4e-07 W=4e-06 AD=1.84e-12 AS=1.4e-13 PD=4.6e-06 PS=2.3e-06 w_cont=6e-07 nfing=1 mmm=1 $X=145240 $Y=155280 $D=5
M1 3 2 1 1 pmos_a L=2.4e-07 W=4e-06 AD=1.84e-12 AS=1.4e-13 PD=4.6e-06 PS=2.3e-06 w_cont=6e-07 nfing=1 mmm=1 $X=159240 $Y=155280 $D=5
M2 3 2 1 1 pmos_a L=2.4e-07 W=4e-06 AD=1.84e-12 AS=1.4e-13 PD=4.6e-06 PS=2.3e-06 w_cont=6e-07 nfing=1 mmm=1 $X=167740 $Y=155280 $D=5
X6 4 1 3 nmos_io_a_CDNS_5887047866531 $T=147560 137260 1 180 $X=144660 $Y=137160
X7 4 1 3 nmos_io_a_CDNS_5887047866531 $T=147560 164660 1 180 $X=144660 $Y=164560
X8 4 1 3 nmos_io_a_CDNS_5887047866531 $T=151660 137260 0 0 $X=151660 $Y=137160
X9 4 1 3 nmos_io_a_CDNS_5887047866531 $T=151660 164660 0 0 $X=151660 $Y=164560
X10 4 1 3 nmos_io_a_CDNS_5887047866531 $T=161560 137260 1 180 $X=158660 $Y=137160
X11 4 1 3 nmos_io_a_CDNS_5887047866531 $T=161560 164660 1 180 $X=158660 $Y=164560
X12 4 1 3 nmos_io_a_CDNS_5887047866531 $T=165660 137260 0 0 $X=165660 $Y=137160
X13 4 1 3 nmos_io_a_CDNS_5887047866531 $T=165660 164660 0 0 $X=165660 $Y=164560
X14 4 3 2 nmos_a_CDNS_5887047866530 $T=151660 155080 0 0 $X=151660 $Y=155080
.ENDS
***************************************
.SUBCKT ICV_60 1 2 3
** N=3 EP=3 IP=12 FDC=4
X0 1 2 3 nmos_io_a_CDNS_5887047866531 $T=147560 109860 1 180 $X=144660 $Y=109760
X1 1 2 3 nmos_io_a_CDNS_5887047866531 $T=151660 109860 0 0 $X=151660 $Y=109760
X2 1 2 3 nmos_io_a_CDNS_5887047866531 $T=161560 109860 1 180 $X=158660 $Y=109760
X3 1 2 3 nmos_io_a_CDNS_5887047866531 $T=165660 109860 0 0 $X=165660 $Y=109760
.ENDS
***************************************
.SUBCKT ICV_61 1 2 3 4
** N=4 EP=4 IP=48 FDC=16
M0 4 2 3 3 pmos_a L=2.4e-07 W=4e-06 AD=1.84e-12 AS=1.4e-13 PD=4.6e-06 PS=2.3e-06 w_cont=6e-07 nfing=1 mmm=1 $X=45280 $Y=-167980 $D=5
M1 4 2 3 3 pmos_a L=2.4e-07 W=4e-06 AD=1.84e-12 AS=1.4e-13 PD=4.6e-06 PS=2.3e-06 w_cont=6e-07 nfing=1 mmm=1 $X=45280 $Y=-159480 $D=5
M2 4 2 3 3 pmos_a L=2.4e-07 W=4e-06 AD=1.84e-12 AS=1.4e-13 PD=4.6e-06 PS=2.3e-06 w_cont=6e-07 nfing=1 mmm=1 $X=45280 $Y=-145480 $D=5
X6 1 3 4 nmos_io_a_CDNS_5887047866531 $T=25660 -165660 0 270 $X=25560 $Y=-168560
X7 1 3 4 nmos_io_a_CDNS_5887047866531 $T=25660 -161560 1 90 $X=25560 $Y=-161560
X8 1 3 4 nmos_io_a_CDNS_5887047866531 $T=25660 -151660 0 270 $X=25560 $Y=-154560
X9 1 3 4 nmos_io_a_CDNS_5887047866531 $T=25660 -147560 1 90 $X=25560 $Y=-147560
X10 1 3 4 nmos_io_a_CDNS_5887047866531 $T=55060 -165660 0 270 $X=54960 $Y=-168560
X11 1 3 4 nmos_io_a_CDNS_5887047866531 $T=55060 -161560 1 90 $X=54960 $Y=-161560
X12 1 3 4 nmos_io_a_CDNS_5887047866531 $T=55060 -151660 0 270 $X=54960 $Y=-154560
X13 1 3 4 nmos_io_a_CDNS_5887047866531 $T=55060 -147560 1 90 $X=54960 $Y=-147560
X14 1 3 4 nmos_io_a_CDNS_5887047866531 $T=82460 -165660 0 270 $X=82360 $Y=-168560
X15 1 3 4 nmos_io_a_CDNS_5887047866531 $T=82460 -161560 1 90 $X=82360 $Y=-161560
X16 1 3 4 nmos_io_a_CDNS_5887047866531 $T=82460 -151660 0 270 $X=82360 $Y=-154560
X17 1 3 4 nmos_io_a_CDNS_5887047866531 $T=82460 -147560 1 90 $X=82360 $Y=-147560
X18 1 4 2 nmos_a_CDNS_5887047866530 $T=43580 -151660 0 270 $X=43580 $Y=-153100
.ENDS
***************************************
.SUBCKT ICV_62 1 2 3
** N=4 EP=3 IP=12 FDC=4
X0 1 2 3 nmos_io_a_CDNS_5887047866531 $T=260 -165660 0 270 $X=160 $Y=-168560
X1 1 2 3 nmos_io_a_CDNS_5887047866531 $T=260 -161560 1 90 $X=160 $Y=-161560
X2 1 2 3 nmos_io_a_CDNS_5887047866531 $T=260 -151660 0 270 $X=160 $Y=-154560
X3 1 2 3 nmos_io_a_CDNS_5887047866531 $T=260 -147560 1 90 $X=160 $Y=-147560
.ENDS
***************************************
.SUBCKT ICV_63 1 2 5
** N=5 EP=3 IP=7 FDC=161
X0 2 1 5 nmos_io_a_CDNS_5887047866531 $T=190400 -137660 0 270 $X=190300 $Y=-140560
X1 1 2 cpoly_n_CDNS_5887047866535 $T=211680 -135500 0 0 $X=211680 $Y=-135500
X2 2 1 cpoly_p_CDNS_5887047866528 $T=211900 -121380 0 0 $X=211900 $Y=-121380
.ENDS
***************************************
.SUBCKT ICV_64 1 2 3 4
** N=4 EP=4 IP=9 FDC=3
M0 4 2 1 1 pmos_a L=2.4e-07 W=4e-06 AD=1.84e-12 AS=1.4e-13 PD=4.6e-06 PS=2.3e-06 w_cont=6e-07 nfing=1 mmm=1 $X=139740 $Y=155280 $D=5
X2 3 1 4 nmos_io_a_CDNS_5887047866531 $T=137660 137260 0 0 $X=137660 $Y=137160
X3 3 1 4 nmos_io_a_CDNS_5887047866531 $T=137660 164660 0 0 $X=137660 $Y=164560
.ENDS
***************************************
.SUBCKT ICV_65 1 2 3 4 5
** N=5 EP=5 IP=33 FDC=11
M0 4 5 2 2 pmos_a L=2.4e-07 W=4e-06 AD=1.84e-12 AS=1.4e-13 PD=4.6e-06 PS=2.3e-06 w_cont=6e-07 nfing=1 mmm=1 $X=118440 $Y=105760 $D=5
M1 4 5 2 2 pmos_a L=2.4e-07 W=4e-06 AD=1.84e-12 AS=1.4e-13 PD=4.6e-06 PS=2.3e-06 w_cont=6e-07 nfing=1 mmm=1 $X=118440 $Y=115000 $D=5
M2 4 5 2 2 pmos_a L=2.4e-07 W=4e-06 AD=1.84e-12 AS=1.4e-13 PD=4.6e-06 PS=2.3e-06 w_cont=6e-07 nfing=1 mmm=1 $X=118440 $Y=124400 $D=5
M3 4 5 2 2 pmos_a L=2.4e-07 W=4e-06 AD=1.84e-12 AS=1.4e-13 PD=4.6e-06 PS=2.3e-06 w_cont=6e-07 nfing=1 mmm=1 $X=118440 $Y=133920 $D=5
M4 4 5 2 2 pmos_a L=2.4e-07 W=4e-06 AD=1.84e-12 AS=1.4e-13 PD=4.6e-06 PS=2.3e-06 w_cont=6e-07 nfing=1 mmm=1 $X=131580 $Y=105760 $D=5
M5 4 5 2 2 pmos_a L=2.4e-07 W=4e-06 AD=1.84e-12 AS=1.4e-13 PD=4.6e-06 PS=2.3e-06 w_cont=6e-07 nfing=1 mmm=1 $X=131580 $Y=115000 $D=5
M6 4 5 2 2 pmos_a L=2.4e-07 W=4e-06 AD=1.84e-12 AS=1.4e-13 PD=4.6e-06 PS=2.3e-06 w_cont=6e-07 nfing=1 mmm=1 $X=131580 $Y=124400 $D=5
M7 4 5 2 2 pmos_a L=2.4e-07 W=4e-06 AD=1.84e-12 AS=1.4e-13 PD=4.6e-06 PS=2.3e-06 w_cont=6e-07 nfing=1 mmm=1 $X=131580 $Y=133920 $D=5
X16 1 2 3 nmos_io_a_CDNS_5887047866531 $T=137660 109860 0 0 $X=137660 $Y=109760
X17 1 4 5 nmos_a_CDNS_5887047866530 $T=119300 94920 1 180 $X=117860 $Y=94920
X18 1 4 5 nmos_a_CDNS_5887047866530 $T=130960 94940 0 0 $X=130960 $Y=94940
.ENDS
***************************************
.SUBCKT ICV_66 1 2 3 4 5
** N=5 EP=5 IP=28 FDC=26
M0 4 3 5 5 pmos_a L=2.4e-07 W=4e-06 AD=1.84e-12 AS=1.4e-13 PD=4.6e-06 PS=2.3e-06 w_cont=6e-07 nfing=1 mmm=1 $X=45280 $Y=-139980 $D=5
X2 1 5 4 nmos_io_a_CDNS_5887047866531 $T=25660 -137660 0 270 $X=25560 $Y=-140560
X3 1 5 4 nmos_io_a_CDNS_5887047866531 $T=55060 -137660 0 270 $X=54960 $Y=-140560
X4 1 5 4 nmos_io_a_CDNS_5887047866531 $T=82460 -137660 0 270 $X=82360 $Y=-140560
X5 1 3 2 nmos_a_CDNS_5887047866530 $T=86980 -130960 0 270 $X=86980 $Y=-132400
X6 1 3 2 nmos_a_CDNS_5887047866530 $T=86980 -119300 1 90 $X=86980 $Y=-119300
X7 2 5 cpoly_p_CDNS_5887047866534 $T=32440 -118720 1 0 $X=32440 $Y=-131220
X8 2 5 cpoly_p_CDNS_5887047866534 $T=43200 -118720 1 0 $X=43200 $Y=-131220
X9 2 5 cpoly_p_CDNS_5887047866534 $T=53960 -118720 1 0 $X=53960 $Y=-131220
X10 2 5 cpoly_p_CDNS_5887047866534 $T=64720 -118720 1 0 $X=64720 $Y=-131220
X11 2 5 cpoly_p_CDNS_5887047866534 $T=75480 -118720 1 0 $X=75480 $Y=-131220
.ENDS
***************************************
.SUBCKT ICV_67 1 2 3 4
** N=5 EP=4 IP=7 FDC=9
X0 1 2 3 nmos_io_a_CDNS_5887047866531 $T=260 -137660 0 270 $X=160 $Y=-140560
X1 4 2 cpoly_p_CDNS_5887047866534 $T=140 -118720 1 0 $X=140 $Y=-131220
X2 4 2 cpoly_p_CDNS_5887047866534 $T=10920 -118720 1 0 $X=10920 $Y=-131220
.ENDS
***************************************
.SUBCKT ICV_68 1 2 5
** N=5 EP=3 IP=11 FDC=83
X0 2 1 5 nmos_io_a_CDNS_5887047866531 $T=190400 -109660 0 270 $X=190300 $Y=-112560
X1 2 1 5 nmos_io_a_CDNS_5887047866531 $T=190400 -105560 1 90 $X=190300 $Y=-105560
X2 2 1 5 nmos_io_a_CDNS_5887047866531 $T=190400 -95660 0 270 $X=190300 $Y=-98560
X3 1 2 cpoly_n_CDNS_5887047866535 $T=211680 -106040 0 0 $X=211680 $Y=-106040
.ENDS
***************************************
.SUBCKT ICV_69 1 2 3 4
** N=4 EP=4 IP=27 FDC=9
M0 4 2 1 1 pmos_a L=2.4e-07 W=4e-06 AD=1.84e-12 AS=1.4e-13 PD=4.6e-06 PS=2.3e-06 w_cont=6e-07 nfing=1 mmm=1 $X=155280 $Y=-111980 $D=5
M1 4 2 1 1 pmos_a L=2.4e-07 W=4e-06 AD=1.84e-12 AS=1.4e-13 PD=4.6e-06 PS=2.3e-06 w_cont=6e-07 nfing=1 mmm=1 $X=155280 $Y=-103480 $D=5
X4 3 1 4 nmos_io_a_CDNS_5887047866531 $T=137260 -109660 0 270 $X=137160 $Y=-112560
X5 3 1 4 nmos_io_a_CDNS_5887047866531 $T=137260 -105560 1 90 $X=137160 $Y=-105560
X6 3 1 4 nmos_io_a_CDNS_5887047866531 $T=137260 -95660 0 270 $X=137160 $Y=-98560
X7 3 1 4 nmos_io_a_CDNS_5887047866531 $T=164660 -109660 0 270 $X=164560 $Y=-112560
X8 3 1 4 nmos_io_a_CDNS_5887047866531 $T=164660 -105560 1 90 $X=164560 $Y=-105560
X9 3 1 4 nmos_io_a_CDNS_5887047866531 $T=164660 -95660 0 270 $X=164560 $Y=-98560
X10 3 4 2 nmos_a_CDNS_5887047866530 $T=155080 -95660 0 270 $X=155080 $Y=-97100
.ENDS
***************************************
.SUBCKT ICV_70 1 2 3
** N=3 EP=3 IP=9 FDC=3
X0 1 2 3 nmos_io_a_CDNS_5887047866531 $T=109860 -109660 0 270 $X=109760 $Y=-112560
X1 1 2 3 nmos_io_a_CDNS_5887047866531 $T=109860 -105560 1 90 $X=109760 $Y=-105560
X2 1 2 3 nmos_io_a_CDNS_5887047866531 $T=109860 -95660 0 270 $X=109760 $Y=-98560
.ENDS
***************************************
.SUBCKT ICV_71 1 2 3 4
** N=4 EP=4 IP=36 FDC=12
M0 4 2 3 3 pmos_a L=2.4e-07 W=4e-06 AD=1.84e-12 AS=1.4e-13 PD=4.6e-06 PS=2.3e-06 w_cont=6e-07 nfing=1 mmm=1 $X=45280 $Y=-111980 $D=5
M1 4 2 3 3 pmos_a L=2.4e-07 W=4e-06 AD=1.84e-12 AS=1.4e-13 PD=4.6e-06 PS=2.3e-06 w_cont=6e-07 nfing=1 mmm=1 $X=45280 $Y=-103480 $D=5
X4 1 3 4 nmos_io_a_CDNS_5887047866531 $T=25720 -109660 0 270 $X=25620 $Y=-112560
X5 1 3 4 nmos_io_a_CDNS_5887047866531 $T=25720 -105560 1 90 $X=25620 $Y=-105560
X6 1 3 4 nmos_io_a_CDNS_5887047866531 $T=25720 -95660 0 270 $X=25620 $Y=-98560
X7 1 3 4 nmos_io_a_CDNS_5887047866531 $T=55060 -109660 0 270 $X=54960 $Y=-112560
X8 1 3 4 nmos_io_a_CDNS_5887047866531 $T=55060 -105560 1 90 $X=54960 $Y=-105560
X9 1 3 4 nmos_io_a_CDNS_5887047866531 $T=55060 -95660 0 270 $X=54960 $Y=-98560
X10 1 3 4 nmos_io_a_CDNS_5887047866531 $T=82460 -109660 0 270 $X=82360 $Y=-112560
X11 1 3 4 nmos_io_a_CDNS_5887047866531 $T=82460 -105560 1 90 $X=82360 $Y=-105560
X12 1 3 4 nmos_io_a_CDNS_5887047866531 $T=82460 -95660 0 270 $X=82360 $Y=-98560
X13 1 4 2 nmos_a_CDNS_5887047866530 $T=43580 -95660 0 270 $X=43580 $Y=-97100
.ENDS
***************************************
.SUBCKT ICV_72 1 2 3
** N=4 EP=3 IP=9 FDC=3
X0 1 2 3 nmos_io_a_CDNS_5887047866531 $T=260 -109660 0 270 $X=160 $Y=-112560
X1 1 2 3 nmos_io_a_CDNS_5887047866531 $T=260 -105560 1 90 $X=160 $Y=-105560
X2 1 2 3 nmos_io_a_CDNS_5887047866531 $T=260 -95660 0 270 $X=160 $Y=-98560
.ENDS
***************************************
.SUBCKT ICV_73 1 2 5
** N=5 EP=3 IP=8 FDC=82
X0 2 1 5 nmos_io_a_CDNS_5887047866531 $T=190400 -91560 1 90 $X=190300 $Y=-91560
X1 2 1 5 nmos_io_a_CDNS_5887047866531 $T=190400 -81660 0 270 $X=190300 $Y=-84560
X2 2 1 cpoly_p_CDNS_5887047866528 $T=211900 -91920 0 0 $X=211900 $Y=-91920
.ENDS
***************************************
.SUBCKT ICV_74 1 2 3 4
** N=4 EP=4 IP=18 FDC=6
M0 4 2 1 1 pmos_a L=2.4e-07 W=4e-06 AD=1.84e-12 AS=1.4e-13 PD=4.6e-06 PS=2.3e-06 w_cont=6e-07 nfing=1 mmm=1 $X=155280 $Y=-89480 $D=5
M1 4 2 1 1 pmos_a L=2.4e-07 W=4e-06 AD=1.84e-12 AS=1.4e-13 PD=4.6e-06 PS=2.3e-06 w_cont=6e-07 nfing=1 mmm=1 $X=155280 $Y=-83980 $D=5
X4 3 1 4 nmos_io_a_CDNS_5887047866531 $T=137260 -91560 1 90 $X=137160 $Y=-91560
X5 3 1 4 nmos_io_a_CDNS_5887047866531 $T=137260 -81660 0 270 $X=137160 $Y=-84560
X6 3 1 4 nmos_io_a_CDNS_5887047866531 $T=164660 -91560 1 90 $X=164560 $Y=-91560
X7 3 1 4 nmos_io_a_CDNS_5887047866531 $T=164660 -81660 0 270 $X=164560 $Y=-84560
.ENDS
***************************************
.SUBCKT ICV_75 1 2 3
** N=3 EP=3 IP=6 FDC=2
X0 1 2 3 nmos_io_a_CDNS_5887047866531 $T=109860 -91560 1 90 $X=109760 $Y=-91560
X1 1 2 3 nmos_io_a_CDNS_5887047866531 $T=109860 -81660 0 270 $X=109760 $Y=-84560
.ENDS
***************************************
.SUBCKT ICV_76 1 2 3 4
** N=4 EP=4 IP=24 FDC=8
M0 3 2 4 4 pmos_a L=2.4e-07 W=4e-06 AD=1.84e-12 AS=1.4e-13 PD=4.6e-06 PS=2.3e-06 w_cont=6e-07 nfing=1 mmm=1 $X=45280 $Y=-89480 $D=5
M1 3 2 4 4 pmos_a L=2.4e-07 W=4e-06 AD=1.84e-12 AS=1.4e-13 PD=4.6e-06 PS=2.3e-06 w_cont=6e-07 nfing=1 mmm=1 $X=45280 $Y=-83980 $D=5
X4 1 4 3 nmos_io_a_CDNS_5887047866531 $T=25720 -91560 1 90 $X=25620 $Y=-91560
X5 1 4 3 nmos_io_a_CDNS_5887047866531 $T=25720 -81660 0 270 $X=25620 $Y=-84560
X6 1 4 3 nmos_io_a_CDNS_5887047866531 $T=55060 -91560 1 90 $X=54960 $Y=-91560
X7 1 4 3 nmos_io_a_CDNS_5887047866531 $T=55060 -81660 0 270 $X=54960 $Y=-84560
X8 1 4 3 nmos_io_a_CDNS_5887047866531 $T=82460 -91560 1 90 $X=82360 $Y=-91560
X9 1 4 3 nmos_io_a_CDNS_5887047866531 $T=82460 -81660 0 270 $X=82360 $Y=-84560
.ENDS
***************************************
.SUBCKT ICV_77 1 2 3
** N=4 EP=3 IP=6 FDC=2
X0 1 2 3 nmos_io_a_CDNS_5887047866531 $T=260 -91560 1 90 $X=160 $Y=-91560
X1 1 2 3 nmos_io_a_CDNS_5887047866531 $T=260 -81660 0 270 $X=160 $Y=-84560
.ENDS
***************************************
.SUBCKT ICV_78
** N=4 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT ICV_79
** N=2 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT ICV_80
** N=2 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT ICV_81
** N=2 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT ICV_82
** N=3 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT PAD_Clamp_200 VDD_PAD vdd! gnd! GND_PAD
** N=8 EP=4 IP=140 FDC=2421
X0 GND_PAD 7 rppoly_CDNS_5887047866532 $T=136620 204240 1 270 $X=132880 $Y=1140
X1 7 VDD_PAD cpoly_p_CDNS_5887047866534 $T=118720 21680 1 90 $X=118720 $Y=21680
X2 vdd! gnd! ICV_40 $T=520 433340 0 0 $X=520 $Y=433340
X3 gnd! vdd! ICV_41 $T=520 420500 0 0 $X=520 $Y=420500
X4 GND_PAD VDD_PAD ICV_42 $T=150840 211900 0 90 $X=142840 $Y=211900
X5 GND_PAD VDD_PAD ICV_43 $T=180440 220 0 90 $X=172440 $Y=220
X6 GND_PAD VDD_PAD ICV_44 $T=67280 220 0 90 $X=59280 $Y=220
X7 GND_PAD VDD_PAD ICV_45 $T=48420 220 0 90 $X=40420 $Y=220
X8 GND_PAD VDD_PAD ICV_46 $T=29560 220 0 90 $X=21560 $Y=220
X9 GND_PAD VDD_PAD ICV_47 $T=10700 220 0 90 $X=2700 $Y=220
X10 GND_PAD VDD_PAD ICV_48 $T=189620 0 0 90 $X=182120 $Y=0
X11 GND_PAD VDD_PAD ICV_49 $T=76460 0 0 90 $X=68960 $Y=0
X12 GND_PAD VDD_PAD ICV_50 $T=57600 0 0 90 $X=50100 $Y=0
X13 GND_PAD VDD_PAD ICV_51 $T=38740 0 0 90 $X=31240 $Y=0
X14 GND_PAD VDD_PAD ICV_52 $T=19880 0 0 90 $X=12380 $Y=0
X20 VDD_PAD GND_PAD 6 ICV_58 $T=0 0 0 90 $X=144660 $Y=179300
X21 VDD_PAD 5 6 GND_PAD ICV_59 $T=0 0 0 0 $X=144620 $Y=137160
X22 GND_PAD VDD_PAD 6 ICV_60 $T=0 0 0 0 $X=144660 $Y=97100
X23 GND_PAD 5 VDD_PAD 6 ICV_61 $T=0 0 0 90 $X=144620 $Y=25560
X24 GND_PAD VDD_PAD 6 ICV_62 $T=0 0 0 90 $X=144660 $Y=-136000
X25 VDD_PAD GND_PAD 6 ICV_63 $T=0 0 0 90 $X=112600 $Y=179300
X26 VDD_PAD 5 GND_PAD 6 ICV_64 $T=0 0 0 0 $X=112600 $Y=137160
X27 GND_PAD VDD_PAD 6 5 7 ICV_65 $T=0 0 0 0 $X=112600 $Y=94920
X28 GND_PAD 7 5 6 VDD_PAD ICV_66 $T=0 0 0 90 $X=112600 $Y=25560
X29 GND_PAD VDD_PAD 6 7 ICV_67 $T=0 0 0 90 $X=112600 $Y=-136000
X30 VDD_PAD GND_PAD 6 ICV_68 $T=0 0 0 90 $X=95660 $Y=179300
X31 VDD_PAD 5 GND_PAD 6 ICV_69 $T=0 0 0 90 $X=95660 $Y=137160
X32 GND_PAD VDD_PAD 6 ICV_70 $T=0 0 0 90 $X=95660 $Y=97100
X33 GND_PAD 5 VDD_PAD 6 ICV_71 $T=0 0 0 90 $X=95660 $Y=25600
X34 GND_PAD VDD_PAD 6 ICV_72 $T=0 0 0 90 $X=95660 $Y=-136000
X35 VDD_PAD GND_PAD 6 ICV_73 $T=0 0 0 90 $X=81660 $Y=179300
X36 VDD_PAD 5 GND_PAD 6 ICV_74 $T=0 0 0 90 $X=81660 $Y=137160
X37 GND_PAD VDD_PAD 6 ICV_75 $T=0 0 0 90 $X=81660 $Y=97100
X38 GND_PAD 5 6 VDD_PAD ICV_76 $T=0 0 0 90 $X=81660 $Y=25600
X39 GND_PAD VDD_PAD 6 ICV_77 $T=0 0 0 90 $X=81660 $Y=-136000
.ENDS
***************************************
.SUBCKT cpoly_p_CDNS_5887047866568 1 2
** N=2 EP=2 IP=0 FDC=1
M0 1 2 1 cpoly_p w=6e-06 l=2e-06 c=8.0712e-14 as=1.68e-13 ad=1.152e-12 ps=1.44e-06 pd=2.27368e-06 sim_w=2.88e-06 m_per_maxw=2.08333 numb_sub_cont=4 nfing=1 $X=620 $Y=200 $D=21
.ENDS
***************************************
.SUBCKT nmos_a_CDNS_5887047866521 1 2 3
** N=3 EP=3 IP=0 FDC=1
M0 2 3 1 1 nmos_a L=2.4e-07 W=5e-07 AD=4.4e-13 AS=2e-13 PD=1.1e-06 PS=5.5e-07 w_cont=6e-07 nfing=1 source_num=2 $X=620 $Y=200 $D=1
.ENDS
***************************************
.SUBCKT cpoly_n_CDNS_5887047866570 1 2
** N=2 EP=2 IP=0 FDC=17
M0 1 2 1 cpoly_n w=6e-06 l=2e-06 c=7.5402e-14 as=2.4e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.4338e-06 sim_w=5.76e-06 m_per_maxw=1.04167 numb_sub_cont=3 nfing=1 $X=620 $Y=200 $D=22
M1 1 2 1 cpoly_n w=6e-06 l=2e-06 c=7.5402e-14 as=3.0336e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.4338e-06 sim_w=5.76e-06 m_per_maxw=1.04167 numb_sub_cont=3 nfing=1 $X=3140 $Y=200 $D=22
M2 1 2 1 cpoly_n w=6e-06 l=2e-06 c=7.5402e-14 as=3.0336e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.4338e-06 sim_w=5.76e-06 m_per_maxw=1.04167 numb_sub_cont=3 nfing=1 $X=5660 $Y=200 $D=22
M3 1 2 1 cpoly_n w=6e-06 l=2e-06 c=7.5402e-14 as=3.0336e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.4338e-06 sim_w=5.76e-06 m_per_maxw=1.04167 numb_sub_cont=3 nfing=1 $X=8180 $Y=200 $D=22
M4 1 2 1 cpoly_n w=6e-06 l=2e-06 c=7.5402e-14 as=3.0336e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.4338e-06 sim_w=5.76e-06 m_per_maxw=1.04167 numb_sub_cont=3 nfing=1 $X=10700 $Y=200 $D=22
M5 1 2 1 cpoly_n w=6e-06 l=2e-06 c=7.5402e-14 as=3.0336e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.4338e-06 sim_w=5.76e-06 m_per_maxw=1.04167 numb_sub_cont=3 nfing=1 $X=13220 $Y=200 $D=22
M6 1 2 1 cpoly_n w=6e-06 l=2e-06 c=7.5402e-14 as=3.0336e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.4338e-06 sim_w=5.76e-06 m_per_maxw=1.04167 numb_sub_cont=3 nfing=1 $X=15740 $Y=200 $D=22
M7 1 2 1 cpoly_n w=6e-06 l=2e-06 c=7.5402e-14 as=3.0336e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.4338e-06 sim_w=5.76e-06 m_per_maxw=1.04167 numb_sub_cont=3 nfing=1 $X=18260 $Y=200 $D=22
M8 1 2 1 cpoly_n w=6e-06 l=2e-06 c=7.5402e-14 as=3.0336e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.4338e-06 sim_w=5.76e-06 m_per_maxw=1.04167 numb_sub_cont=3 nfing=1 $X=20780 $Y=200 $D=22
M9 1 2 1 cpoly_n w=6e-06 l=2e-06 c=7.5402e-14 as=3.0336e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.4338e-06 sim_w=5.76e-06 m_per_maxw=1.04167 numb_sub_cont=3 nfing=1 $X=23300 $Y=200 $D=22
M10 1 2 1 cpoly_n w=6e-06 l=2e-06 c=7.5402e-14 as=3.0336e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.4338e-06 sim_w=5.76e-06 m_per_maxw=1.04167 numb_sub_cont=3 nfing=1 $X=25820 $Y=200 $D=22
M11 1 2 1 cpoly_n w=6e-06 l=2e-06 c=7.5402e-14 as=3.0336e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.4338e-06 sim_w=5.76e-06 m_per_maxw=1.04167 numb_sub_cont=3 nfing=1 $X=28340 $Y=200 $D=22
M12 1 2 1 cpoly_n w=6e-06 l=2e-06 c=7.5402e-14 as=3.0336e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.4338e-06 sim_w=5.76e-06 m_per_maxw=1.04167 numb_sub_cont=3 nfing=1 $X=30860 $Y=200 $D=22
M13 1 2 1 cpoly_n w=6e-06 l=2e-06 c=7.5402e-14 as=3.0336e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.4338e-06 sim_w=5.76e-06 m_per_maxw=1.04167 numb_sub_cont=3 nfing=1 $X=33380 $Y=200 $D=22
M14 1 2 1 cpoly_n w=6e-06 l=2e-06 c=7.5402e-14 as=3.0336e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.4338e-06 sim_w=5.76e-06 m_per_maxw=1.04167 numb_sub_cont=3 nfing=1 $X=35900 $Y=200 $D=22
M15 1 2 1 cpoly_n w=6e-06 l=2e-06 c=7.5402e-14 as=3.0336e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.4338e-06 sim_w=5.76e-06 m_per_maxw=1.04167 numb_sub_cont=3 nfing=1 $X=38420 $Y=200 $D=22
M16 1 2 1 cpoly_n w=6e-06 l=2e-06 c=7.5402e-14 as=3.0336e-13 ad=2.304e-12 ps=2.88e-06 pd=4.86761e-06 sim_w=5.76e-06 m_per_maxw=1.04167 numb_sub_cont=3 nfing=1 $X=40940 $Y=200 $D=22
.ENDS
***************************************
.SUBCKT cpoly_p_CDNS_5887047866569 1 2
** N=2 EP=2 IP=0 FDC=17
M0 1 2 1 cpoly_p w=6e-06 l=2e-06 c=8.0712e-14 as=1.68e-13 ad=7.488e-13 ps=1.44e-06 pd=1.13684e-06 sim_w=2.88e-06 m_per_maxw=2.08333 numb_sub_cont=4 nfing=1 $X=620 $Y=200 $D=21
M1 1 2 1 cpoly_p w=6e-06 l=2e-06 c=8.0712e-14 as=2.1408e-13 ad=7.488e-13 ps=1.44e-06 pd=1.13684e-06 sim_w=2.88e-06 m_per_maxw=2.08333 numb_sub_cont=4 nfing=1 $X=3140 $Y=200 $D=21
M2 1 2 1 cpoly_p w=6e-06 l=2e-06 c=8.0712e-14 as=2.1408e-13 ad=7.488e-13 ps=1.44e-06 pd=1.13684e-06 sim_w=2.88e-06 m_per_maxw=2.08333 numb_sub_cont=4 nfing=1 $X=5660 $Y=200 $D=21
M3 1 2 1 cpoly_p w=6e-06 l=2e-06 c=8.0712e-14 as=2.1408e-13 ad=7.488e-13 ps=1.44e-06 pd=1.13684e-06 sim_w=2.88e-06 m_per_maxw=2.08333 numb_sub_cont=4 nfing=1 $X=8180 $Y=200 $D=21
M4 1 2 1 cpoly_p w=6e-06 l=2e-06 c=8.0712e-14 as=2.1408e-13 ad=7.488e-13 ps=1.44e-06 pd=1.13684e-06 sim_w=2.88e-06 m_per_maxw=2.08333 numb_sub_cont=4 nfing=1 $X=10700 $Y=200 $D=21
M5 1 2 1 cpoly_p w=6e-06 l=2e-06 c=8.0712e-14 as=2.1408e-13 ad=7.488e-13 ps=1.44e-06 pd=1.13684e-06 sim_w=2.88e-06 m_per_maxw=2.08333 numb_sub_cont=4 nfing=1 $X=13220 $Y=200 $D=21
M6 1 2 1 cpoly_p w=6e-06 l=2e-06 c=8.0712e-14 as=2.1408e-13 ad=7.488e-13 ps=1.44e-06 pd=1.13684e-06 sim_w=2.88e-06 m_per_maxw=2.08333 numb_sub_cont=4 nfing=1 $X=15740 $Y=200 $D=21
M7 1 2 1 cpoly_p w=6e-06 l=2e-06 c=8.0712e-14 as=2.1408e-13 ad=7.488e-13 ps=1.44e-06 pd=1.13684e-06 sim_w=2.88e-06 m_per_maxw=2.08333 numb_sub_cont=4 nfing=1 $X=18260 $Y=200 $D=21
M8 1 2 1 cpoly_p w=6e-06 l=2e-06 c=8.0712e-14 as=2.1408e-13 ad=7.488e-13 ps=1.44e-06 pd=1.13684e-06 sim_w=2.88e-06 m_per_maxw=2.08333 numb_sub_cont=4 nfing=1 $X=20780 $Y=200 $D=21
M9 1 2 1 cpoly_p w=6e-06 l=2e-06 c=8.0712e-14 as=2.1408e-13 ad=7.488e-13 ps=1.44e-06 pd=1.13684e-06 sim_w=2.88e-06 m_per_maxw=2.08333 numb_sub_cont=4 nfing=1 $X=23300 $Y=200 $D=21
M10 1 2 1 cpoly_p w=6e-06 l=2e-06 c=8.0712e-14 as=2.1408e-13 ad=7.488e-13 ps=1.44e-06 pd=1.13684e-06 sim_w=2.88e-06 m_per_maxw=2.08333 numb_sub_cont=4 nfing=1 $X=25820 $Y=200 $D=21
M11 1 2 1 cpoly_p w=6e-06 l=2e-06 c=8.0712e-14 as=2.1408e-13 ad=7.488e-13 ps=1.44e-06 pd=1.13684e-06 sim_w=2.88e-06 m_per_maxw=2.08333 numb_sub_cont=4 nfing=1 $X=28340 $Y=200 $D=21
M12 1 2 1 cpoly_p w=6e-06 l=2e-06 c=8.0712e-14 as=2.1408e-13 ad=7.488e-13 ps=1.44e-06 pd=1.13684e-06 sim_w=2.88e-06 m_per_maxw=2.08333 numb_sub_cont=4 nfing=1 $X=30860 $Y=200 $D=21
M13 1 2 1 cpoly_p w=6e-06 l=2e-06 c=8.0712e-14 as=2.1408e-13 ad=7.488e-13 ps=1.44e-06 pd=1.13684e-06 sim_w=2.88e-06 m_per_maxw=2.08333 numb_sub_cont=4 nfing=1 $X=33380 $Y=200 $D=21
M14 1 2 1 cpoly_p w=6e-06 l=2e-06 c=8.0712e-14 as=2.1408e-13 ad=7.488e-13 ps=1.44e-06 pd=1.13684e-06 sim_w=2.88e-06 m_per_maxw=2.08333 numb_sub_cont=4 nfing=1 $X=35900 $Y=200 $D=21
M15 1 2 1 cpoly_p w=6e-06 l=2e-06 c=8.0712e-14 as=2.1408e-13 ad=7.488e-13 ps=1.44e-06 pd=1.13684e-06 sim_w=2.88e-06 m_per_maxw=2.08333 numb_sub_cont=4 nfing=1 $X=38420 $Y=200 $D=21
M16 1 2 1 cpoly_p w=6e-06 l=2e-06 c=8.0712e-14 as=2.1408e-13 ad=1.152e-12 ps=1.44e-06 pd=2.27368e-06 sim_w=2.88e-06 m_per_maxw=2.08333 numb_sub_cont=4 nfing=1 $X=40940 $Y=200 $D=21
.ENDS
***************************************
.SUBCKT cpoly_n_CDNS_5887047866571 1 2
** N=2 EP=2 IP=0 FDC=2
M0 1 2 1 cpoly_n w=6e-06 l=2e-06 c=7.5402e-14 as=2.4e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.4338e-06 sim_w=5.76e-06 m_per_maxw=1.04167 numb_sub_cont=3 nfing=1 $X=620 $Y=200 $D=22
M1 1 2 1 cpoly_n w=6e-06 l=2e-06 c=7.5402e-14 as=2.4e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.4338e-06 sim_w=5.76e-06 m_per_maxw=1.04167 numb_sub_cont=3 nfing=1 $X=3140 $Y=200 $D=22
.ENDS
***************************************
.SUBCKT PADIN_Adress_Select nClk gnd! vdd! A nATD nSelect2 nSelect1 Adr
** N=30 EP=8 IP=191 FDC=205
M0 nATD 22 gnd! gnd! nmos_a L=2.4e-07 W=3.6e-06 AD=1.664e-12 AS=1.44e-12 PD=4.16e-06 PS=2.08e-06 w_cont=1.6e-06 nfing=1 source_num=2 $X=15140 $Y=324580 $D=1
M1 Adr 16 gnd! gnd! nmos_a L=2.4e-07 W=7.2e-06 AD=1.648e-12 AS=2.88e-12 PD=4.12e-06 PS=2.06e-06 w_cont=3.1e-06 nfing=1 source_num=2 $X=60100 $Y=319220 $D=1
M2 Adr 16 gnd! gnd! nmos_a L=2.4e-07 W=7.2e-06 AD=1.648e-12 AS=2.88e-12 PD=4.12e-06 PS=2.06e-06 w_cont=3.1e-06 nfing=1 source_num=2 $X=64840 $Y=319220 $D=1
M3 Adr 16 gnd! gnd! nmos_a L=2.4e-07 W=7.2e-06 AD=1.648e-12 AS=2.88e-12 PD=4.12e-06 PS=2.06e-06 w_cont=3.1e-06 nfing=1 source_num=2 $X=69740 $Y=319220 $D=1
M4 Adr 16 gnd! gnd! nmos_a L=2.4e-07 W=7.2e-06 AD=1.648e-12 AS=2.88e-12 PD=4.12e-06 PS=2.06e-06 w_cont=3.1e-06 nfing=1 source_num=2 $X=74480 $Y=319220 $D=1
M5 Adr 16 gnd! gnd! nmos_a L=2.4e-07 W=7.2e-06 AD=1.648e-12 AS=2.88e-12 PD=4.12e-06 PS=2.06e-06 w_cont=3.1e-06 nfing=1 source_num=2 $X=79380 $Y=319220 $D=1
M6 Adr 16 gnd! gnd! nmos_a L=2.4e-07 W=7.2e-06 AD=1.648e-12 AS=2.88e-12 PD=4.12e-06 PS=2.06e-06 w_cont=3.1e-06 nfing=1 source_num=2 $X=84120 $Y=319220 $D=1
M7 Adr 16 gnd! gnd! nmos_a L=2.4e-07 W=7.2e-06 AD=1.648e-12 AS=2.88e-12 PD=4.12e-06 PS=2.06e-06 w_cont=3.1e-06 nfing=1 source_num=2 $X=89020 $Y=319220 $D=1
M8 Adr 16 gnd! gnd! nmos_a L=2.4e-07 W=7.2e-06 AD=1.648e-12 AS=2.88e-12 PD=4.12e-06 PS=2.06e-06 w_cont=3.1e-06 nfing=1 source_num=2 $X=93760 $Y=319220 $D=1
M9 26 11 gnd! gnd! nmos_a L=2.4e-07 W=2.4e-06 AD=1.4e-12 AS=9.6e-13 PD=3.5e-06 PS=1.75e-06 w_cont=1.1e-06 nfing=1 source_num=2 $X=33840 $Y=326820 $D=1
M10 15 13 26 26 nmos_a L=2.4e-07 W=2.4e-06 AD=1.4e-12 AS=9.6e-13 PD=3.5e-06 PS=1.75e-06 w_cont=1.1e-06 nfing=1 source_num=2 $X=35280 $Y=326540 $D=1
M11 11 30 gnd! gnd! nmos_a L=2.4e-07 W=1.2e-06 AD=7.2e-13 AS=4.8e-13 PD=1.8e-06 PS=9e-07 w_cont=6e-07 nfing=1 source_num=2 $X=9380 $Y=325780 $D=1
M12 18 12 gnd! gnd! nmos_a L=2.4e-07 W=1.2e-06 AD=7.2e-13 AS=4.8e-13 PD=1.8e-06 PS=9e-07 w_cont=6e-07 nfing=1 source_num=2 $X=10820 $Y=325780 $D=1
M13 10 11 18 18 nmos_a L=2.4e-07 W=1.2e-06 AD=4.68e-13 AS=4.8e-13 PD=9e-07 PS=9e-07 w_cont=6e-07 nfing=1 source_num=2 $X=12320 $Y=328520 $D=1
M14 10 9 21 21 nmos_a L=2.4e-07 W=1.2e-06 AD=4.68e-13 AS=4.8e-13 PD=9e-07 PS=9e-07 w_cont=6e-07 nfing=1 source_num=2 $X=13080 $Y=328520 $D=1
M15 21 15 gnd! gnd! nmos_a L=2.4e-07 W=1.2e-06 AD=7.2e-13 AS=4.8e-13 PD=1.8e-06 PS=9e-07 w_cont=6e-07 nfing=1 source_num=2 $X=13700 $Y=325780 $D=1
M16 22 23 gnd! gnd! nmos_a L=2.4e-07 W=1.2e-06 AD=7.2e-13 AS=4.8e-13 PD=1.8e-06 PS=9e-07 w_cont=6e-07 nfing=1 source_num=2 $X=16540 $Y=327840 $D=1
M17 10 25 22 22 nmos_a L=2.4e-07 W=1.2e-06 AD=7.2e-13 AS=4.8e-13 PD=1.8e-06 PS=9e-07 w_cont=6e-07 nfing=1 source_num=2 $X=17980 $Y=331060 $D=1
M18 23 25 gnd! gnd! nmos_a L=2.4e-07 W=1.2e-06 AD=7.2e-13 AS=4.8e-13 PD=1.8e-06 PS=9e-07 w_cont=6e-07 nfing=1 source_num=2 $X=19420 $Y=327840 $D=1
M19 12 15 gnd! gnd! nmos_a L=2.4e-07 W=1.2e-06 AD=7.2e-13 AS=6.24e-13 PD=1.8e-06 PS=9e-07 w_cont=6e-07 nfing=1 source_num=2 $X=36680 $Y=327740 $D=1
M20 28 12 gnd! gnd! nmos_a L=2.4e-07 W=1.2e-06 AD=7.2e-13 AS=6.24e-13 PD=1.8e-06 PS=9e-07 w_cont=6e-07 nfing=1 source_num=2 $X=37440 $Y=327740 $D=1
M21 15 14 28 28 nmos_a L=2.4e-07 W=1.2e-06 AD=7.2e-13 AS=4.8e-13 PD=1.8e-06 PS=9e-07 w_cont=6e-07 nfing=1 source_num=2 $X=38880 $Y=327420 $D=1
M22 13 14 gnd! gnd! nmos_a L=2.4e-07 W=1.2e-06 AD=7.2e-13 AS=4.8e-13 PD=1.8e-06 PS=9e-07 w_cont=6e-07 nfing=1 source_num=2 $X=40280 $Y=327420 $D=1
M23 14 nClk gnd! gnd! nmos_a L=2.4e-07 W=1.2e-06 AD=7.2e-13 AS=4.8e-13 PD=1.8e-06 PS=9e-07 w_cont=6e-07 nfing=1 source_num=2 $X=41720 $Y=327420 $D=1
M24 9 11 gnd! gnd! nmos_a L=2.4e-07 W=4.8e-07 AD=4.32e-13 AS=1.92e-13 PD=1.08e-06 PS=5.4e-07 w_cont=6e-07 nfing=1 source_num=2 $X=12260 $Y=325980 $D=1
M25 16 15 gnd! gnd! nmos_a L=2.4e-07 W=3.6e-06 AD=1.664e-12 AS=1.44e-12 PD=4.16e-06 PS=2.08e-06 w_cont=1.6e-06 nfing=1 source_num=2 $X=47800 $Y=327560 $D=1
M26 16 15 gnd! gnd! nmos_a L=2.4e-07 W=3.6e-06 AD=1.664e-12 AS=1.44e-12 PD=4.16e-06 PS=2.08e-06 w_cont=1.6e-06 nfing=1 source_num=2 $X=53880 $Y=327560 $D=1
M27 20 12 vdd! vdd! pmos_a L=2.4e-07 W=2e-06 AD=1.04e-12 AS=1.3e-13 PD=2.6e-06 PS=1.3e-06 w_cont=6e-07 nfing=1 mmm=1 $X=13640 $Y=334500 $D=5
M28 nATD 22 vdd! vdd! pmos_a L=2.4e-07 W=5.76e-06 AD=2.744e-12 AS=2.488e-13 PD=6.86e-06 PS=3.43e-06 w_cont=1.1e-06 nfing=1 mmm=1 $X=15140 $Y=330600 $D=5
M29 Adr 16 vdd! vdd! pmos_a L=2.4e-07 W=1.1e-05 AD=2.63913e-12 AS=1.96364e-13 PD=6.59782e-06 PS=3.29891e-06 w_cont=1.6e-06 nfing=1 mmm=1 $X=60100 $Y=330700 $D=5
M30 Adr 16 vdd! vdd! pmos_a L=2.4e-07 W=1.1e-05 AD=2.63913e-12 AS=1.96364e-13 PD=6.59782e-06 PS=3.29891e-06 w_cont=1.6e-06 nfing=1 mmm=1 $X=64840 $Y=330700 $D=5
M31 Adr 16 vdd! vdd! pmos_a L=2.4e-07 W=1.1e-05 AD=2.63913e-12 AS=1.96364e-13 PD=6.59782e-06 PS=3.29891e-06 w_cont=1.6e-06 nfing=1 mmm=1 $X=69740 $Y=330700 $D=5
M32 Adr 16 vdd! vdd! pmos_a L=2.4e-07 W=1.088e-05 AD=2.64282e-12 AS=1.98212e-13 PD=6.60706e-06 PS=3.30353e-06 w_cont=1.6e-06 nfing=1 mmm=1 $X=74480 $Y=330820 $D=5
M33 Adr 16 vdd! vdd! pmos_a L=2.4e-07 W=1.1e-05 AD=2.63913e-12 AS=1.96364e-13 PD=6.59782e-06 PS=3.29891e-06 w_cont=1.6e-06 nfing=1 mmm=1 $X=79380 $Y=330700 $D=5
M34 Adr 16 vdd! vdd! pmos_a L=2.4e-07 W=1.1e-05 AD=2.63913e-12 AS=1.96364e-13 PD=6.59782e-06 PS=3.29891e-06 w_cont=1.6e-06 nfing=1 mmm=1 $X=84120 $Y=330700 $D=5
M35 Adr 16 vdd! vdd! pmos_a L=2.4e-07 W=1.1e-05 AD=2.63913e-12 AS=1.96364e-13 PD=6.59782e-06 PS=3.29891e-06 w_cont=1.6e-06 nfing=1 mmm=1 $X=89020 $Y=330700 $D=5
M36 Adr 16 vdd! vdd! pmos_a L=2.4e-07 W=1.1e-05 AD=2.63913e-12 AS=1.96364e-13 PD=6.59782e-06 PS=3.29891e-06 w_cont=1.6e-06 nfing=1 mmm=1 $X=93760 $Y=330700 $D=5
M37 16 15 vdd! vdd! pmos_a L=2.4e-07 W=5.76e-06 AD=2.744e-12 AS=2.488e-13 PD=6.86e-06 PS=3.43e-06 w_cont=1.1e-06 nfing=1 mmm=1 $X=46400 $Y=327560 $D=5
M38 16 15 vdd! vdd! pmos_a L=2.4e-07 W=5.76e-06 AD=2.744e-12 AS=2.488e-13 PD=6.86e-06 PS=3.43e-06 w_cont=1.1e-06 nfing=1 mmm=1 $X=52480 $Y=327560 $D=5
M39 17 17 vdd! vdd! pmos_a L=2.4e-07 W=2e-06 AD=6.76e-13 AS=1.3e-13 PD=1.3e-06 PS=1.3e-06 w_cont=6e-07 nfing=1 mmm=1 $X=9240 $Y=334300 $D=5
M40 17 17 vdd! vdd! pmos_a L=2.4e-07 W=2e-06 AD=6.76e-13 AS=1.66e-13 PD=1.3e-06 PS=1.3e-06 w_cont=6e-07 nfing=1 mmm=1 $X=10000 $Y=334300 $D=5
M41 19 15 vdd! vdd! pmos_a L=2.4e-07 W=2e-06 AD=1.04e-12 AS=1.66e-13 PD=2.6e-06 PS=1.3e-06 w_cont=6e-07 nfing=1 mmm=1 $X=10760 $Y=334300 $D=5
M42 10 11 19 19 pmos_a L=2.4e-07 W=2e-06 AD=6.76e-13 AS=1.3e-13 PD=1.3e-06 PS=1.3e-06 w_cont=6e-07 nfing=1 mmm=1 $X=12320 $Y=331000 $D=5
M43 10 9 20 20 pmos_a L=2.4e-07 W=2e-06 AD=6.76e-13 AS=1.3e-13 PD=1.3e-06 PS=1.3e-06 w_cont=6e-07 nfing=1 mmm=1 $X=13080 $Y=331000 $D=5
M44 22 23 10 10 pmos_a L=2.4e-07 W=2e-06 AD=1.04e-12 AS=1.3e-13 PD=2.6e-06 PS=1.3e-06 w_cont=6e-07 nfing=1 mmm=1 $X=16540 $Y=330600 $D=5
M45 23 25 vdd! vdd! pmos_a L=2.4e-07 W=2e-06 AD=1.04e-12 AS=1.3e-13 PD=2.6e-06 PS=1.3e-06 w_cont=6e-07 nfing=1 mmm=1 $X=19420 $Y=331060 $D=5
M46 25 nSelect2 24 24 pmos_a L=2.4e-07 W=2e-06 AD=1.04e-12 AS=1.3e-13 PD=2.6e-06 PS=1.3e-06 w_cont=6e-07 nfing=1 mmm=1 $X=20860 $Y=331560 $D=5
M47 24 nSelect1 vdd! vdd! pmos_a L=2.4e-07 W=2e-06 AD=1.04e-12 AS=1.3e-13 PD=2.6e-06 PS=1.3e-06 w_cont=6e-07 nfing=1 mmm=1 $X=22300 $Y=331560 $D=5
M48 12 15 vdd! vdd! pmos_a L=2.4e-07 W=2e-06 AD=1.04e-12 AS=1.66e-13 PD=2.6e-06 PS=1.3e-06 w_cont=6e-07 nfing=1 mmm=1 $X=36680 $Y=330700 $D=5
M49 29 12 vdd! vdd! pmos_a L=2.4e-07 W=2e-06 AD=1.04e-12 AS=1.66e-13 PD=2.6e-06 PS=1.3e-06 w_cont=6e-07 nfing=1 mmm=1 $X=37440 $Y=330700 $D=5
M50 15 13 29 29 pmos_a L=2.4e-07 W=2e-06 AD=1.04e-12 AS=1.3e-13 PD=2.6e-06 PS=1.3e-06 w_cont=6e-07 nfing=1 mmm=1 $X=38880 $Y=330200 $D=5
M51 13 14 vdd! vdd! pmos_a L=2.4e-07 W=2e-06 AD=1.04e-12 AS=1.3e-13 PD=2.6e-06 PS=1.3e-06 w_cont=6e-07 nfing=1 mmm=1 $X=40280 $Y=330200 $D=5
M52 14 nClk vdd! vdd! pmos_a L=2.4e-07 W=2e-06 AD=1.04e-12 AS=1.3e-13 PD=2.6e-06 PS=1.3e-06 w_cont=6e-07 nfing=1 mmm=1 $X=41720 $Y=331700 $D=5
M53 9 11 vdd! vdd! pmos_a L=2.4e-07 W=1e-06 AD=6.4e-13 AS=1.25e-13 PD=1.6e-06 PS=8e-07 w_cont=6e-07 nfing=1 mmm=1 $X=12200 $Y=335000 $D=5
M54 17 9 vdd! vdd! pmos_a L=2.4e-07 W=4e-06 AD=1.84e-12 AS=1.4e-13 PD=4.6e-06 PS=2.3e-06 w_cont=6e-07 nfing=1 mmm=1 $X=8800 $Y=329000 $D=5
M55 11 30 17 17 pmos_a L=2.4e-07 W=4e-06 AD=1.84e-12 AS=1.4e-13 PD=4.6e-06 PS=2.3e-06 w_cont=6e-07 nfing=1 mmm=1 $X=10240 $Y=328320 $D=5
M56 27 11 vdd! vdd! pmos_a L=2.4e-07 W=4e-06 AD=1.84e-12 AS=1.4e-13 PD=4.6e-06 PS=2.3e-06 w_cont=6e-07 nfing=1 mmm=1 $X=33840 $Y=331020 $D=5
M57 15 14 27 27 pmos_a L=2.4e-07 W=4e-06 AD=1.84e-12 AS=1.4e-13 PD=4.6e-06 PS=2.3e-06 w_cont=6e-07 nfing=1 mmm=1 $X=35280 $Y=331020 $D=5
M58 vdd! gnd! vdd! cpoly_n w=6e-06 l=2e-06 c=7.5402e-14 as=2.4e-13 ad=2.304e-12 ps=2.88e-06 pd=4.86761e-06 sim_w=5.76e-06 m_per_maxw=1.04167 numb_sub_cont=3 nfing=1 $X=30600 $Y=328520 $D=22
M59 vdd! gnd! vdd! cpoly_n w=6e-06 l=2e-06 c=7.5402e-14 as=2.4e-13 ad=2.304e-12 ps=2.88e-06 pd=4.86761e-06 sim_w=5.76e-06 m_per_maxw=1.04167 numb_sub_cont=3 nfing=1 $X=43200 $Y=328200 $D=22
M60 vdd! gnd! vdd! cpoly_n w=6e-06 l=2e-06 c=7.5402e-14 as=2.4e-13 ad=2.304e-12 ps=2.88e-06 pd=4.86761e-06 sim_w=5.76e-06 m_per_maxw=1.04167 numb_sub_cont=3 nfing=1 $X=49280 $Y=328200 $D=22
M61 vdd! gnd! vdd! cpoly_n w=6e-06 l=2e-06 c=7.5402e-14 as=2.4e-13 ad=2.304e-12 ps=2.88e-06 pd=4.86761e-06 sim_w=5.76e-06 m_per_maxw=1.04167 numb_sub_cont=3 nfing=1 $X=55360 $Y=328200 $D=22
M62 vdd! gnd! vdd! cpoly_n w=6e-06 l=2e-06 c=7.5402e-14 as=2.4e-13 ad=2.304e-12 ps=2.88e-06 pd=4.86761e-06 sim_w=5.76e-06 m_per_maxw=1.04167 numb_sub_cont=3 nfing=1 $X=61600 $Y=328200 $D=22
M63 vdd! gnd! vdd! cpoly_n w=6e-06 l=2e-06 c=7.5402e-14 as=2.4e-13 ad=2.304e-12 ps=2.88e-06 pd=4.86761e-06 sim_w=5.76e-06 m_per_maxw=1.04167 numb_sub_cont=3 nfing=1 $X=61600 $Y=336700 $D=22
M64 vdd! gnd! vdd! cpoly_n w=6e-06 l=2e-06 c=7.5402e-14 as=2.4e-13 ad=2.304e-12 ps=2.88e-06 pd=4.86761e-06 sim_w=5.76e-06 m_per_maxw=1.04167 numb_sub_cont=3 nfing=1 $X=66480 $Y=336700 $D=22
M65 vdd! gnd! vdd! cpoly_n w=6e-06 l=2e-06 c=7.5402e-14 as=2.4e-13 ad=2.304e-12 ps=2.88e-06 pd=4.86761e-06 sim_w=5.76e-06 m_per_maxw=1.04167 numb_sub_cont=3 nfing=1 $X=71240 $Y=328200 $D=22
M66 vdd! gnd! vdd! cpoly_n w=6e-06 l=2e-06 c=7.5402e-14 as=2.4e-13 ad=2.304e-12 ps=2.88e-06 pd=4.86761e-06 sim_w=5.76e-06 m_per_maxw=1.04167 numb_sub_cont=3 nfing=1 $X=71240 $Y=336700 $D=22
M67 vdd! gnd! vdd! cpoly_n w=6e-06 l=2e-06 c=7.5402e-14 as=2.4e-13 ad=2.304e-12 ps=2.88e-06 pd=4.86761e-06 sim_w=5.76e-06 m_per_maxw=1.04167 numb_sub_cont=3 nfing=1 $X=76120 $Y=336700 $D=22
M68 vdd! gnd! vdd! cpoly_n w=6e-06 l=2e-06 c=7.5402e-14 as=2.4e-13 ad=2.304e-12 ps=2.88e-06 pd=4.86761e-06 sim_w=5.76e-06 m_per_maxw=1.04167 numb_sub_cont=3 nfing=1 $X=80880 $Y=328200 $D=22
M69 vdd! gnd! vdd! cpoly_n w=6e-06 l=2e-06 c=7.5402e-14 as=2.4e-13 ad=2.304e-12 ps=2.88e-06 pd=4.86761e-06 sim_w=5.76e-06 m_per_maxw=1.04167 numb_sub_cont=3 nfing=1 $X=80880 $Y=336700 $D=22
M70 vdd! gnd! vdd! cpoly_n w=6e-06 l=2e-06 c=7.5402e-14 as=2.4e-13 ad=2.304e-12 ps=2.88e-06 pd=4.86761e-06 sim_w=5.76e-06 m_per_maxw=1.04167 numb_sub_cont=3 nfing=1 $X=85760 $Y=336700 $D=22
M71 vdd! gnd! vdd! cpoly_n w=6e-06 l=2e-06 c=7.5402e-14 as=2.4e-13 ad=2.304e-12 ps=2.88e-06 pd=4.86761e-06 sim_w=5.76e-06 m_per_maxw=1.04167 numb_sub_cont=3 nfing=1 $X=90520 $Y=328200 $D=22
M72 vdd! gnd! vdd! cpoly_n w=6e-06 l=2e-06 c=7.5402e-14 as=2.4e-13 ad=2.304e-12 ps=2.88e-06 pd=4.86761e-06 sim_w=5.76e-06 m_per_maxw=1.04167 numb_sub_cont=3 nfing=1 $X=90520 $Y=336700 $D=22
M73 vdd! gnd! vdd! cpoly_n w=6e-06 l=2e-06 c=7.5402e-14 as=2.4e-13 ad=2.304e-12 ps=2.88e-06 pd=4.86761e-06 sim_w=5.76e-06 m_per_maxw=1.04167 numb_sub_cont=3 nfing=1 $X=95400 $Y=336700 $D=22
D74 A vdd! dn PJ=0.0002 m=1 $X=4020 $Y=-95300 $D=8
D75 A vdd! dn PJ=0.0002 m=1 $X=4020 $Y=114700 $D=8
D76 gnd! A dn PJ=0.0002 m=1 $X=6340 $Y=-99700 $D=8
D77 gnd! A dn PJ=0.0002 m=1 $X=6340 $Y=110300 $D=8
D78 A vdd! dn PJ=0.0002 m=1 $X=8660 $Y=-95300 $D=8
D79 A vdd! dn PJ=0.0002 m=1 $X=8660 $Y=114700 $D=8
D80 gnd! A dn PJ=0.0001 m=1 $X=10980 $Y=-99700 $D=8
D81 gnd! A dn PJ=0.0001 m=1 $X=10980 $Y=110300 $D=8
D82 A vdd! dn PJ=0.0001 m=1 $X=14160 $Y=4700 $D=8
D83 A vdd! dn PJ=0.0001 m=1 $X=14160 $Y=214700 $D=8
D84 gnd! A dn PJ=0.0002 m=1 $X=16480 $Y=-99700 $D=8
D85 gnd! A dn PJ=0.0002 m=1 $X=16480 $Y=110300 $D=8
D86 A vdd! dn PJ=0.0002 m=1 $X=18800 $Y=-95300 $D=8
D87 A vdd! dn PJ=0.0002 m=1 $X=18800 $Y=114700 $D=8
D88 gnd! A dn PJ=0.0002 m=1 $X=21120 $Y=-99700 $D=8
D89 gnd! A dn PJ=0.0002 m=1 $X=21120 $Y=110300 $D=8
D90 A vdd! dn PJ=0.0002 m=1 $X=23440 $Y=-95300 $D=8
D91 A vdd! dn PJ=0.0002 m=1 $X=23440 $Y=114700 $D=8
D92 gnd! A dn PJ=0.0001 m=1 $X=25760 $Y=-99700 $D=8
D93 gnd! A dn PJ=0.0001 m=1 $X=25760 $Y=110300 $D=8
D94 A vdd! dn PJ=0.0001 m=1 $X=28940 $Y=4700 $D=8
D95 A vdd! dn PJ=0.0001 m=1 $X=28940 $Y=214700 $D=8
D96 gnd! A dn PJ=0.0002 m=1 $X=31260 $Y=-99700 $D=8
D97 gnd! A dn PJ=0.0002 m=1 $X=31260 $Y=110300 $D=8
D98 A vdd! dn PJ=0.0002 m=1 $X=33580 $Y=-95300 $D=8
D99 A vdd! dn PJ=0.0002 m=1 $X=33580 $Y=114700 $D=8
D100 gnd! A dn PJ=0.0002 m=1 $X=35900 $Y=-99700 $D=8
D101 gnd! A dn PJ=0.0002 m=1 $X=35900 $Y=110300 $D=8
D102 A vdd! dn PJ=0.0002 m=1 $X=38220 $Y=-95300 $D=8
D103 A vdd! dn PJ=0.0002 m=1 $X=38220 $Y=114700 $D=8
D104 gnd! A dn PJ=0.0001 m=1 $X=40540 $Y=-99700 $D=8
D105 gnd! A dn PJ=0.0001 m=1 $X=40540 $Y=110300 $D=8
D106 A vdd! dn PJ=0.0001 m=1 $X=43720 $Y=4700 $D=8
D107 A vdd! dn PJ=0.0001 m=1 $X=43720 $Y=214700 $D=8
D108 gnd! A dn PJ=0.0002 m=1 $X=46040 $Y=-99700 $D=8
D109 gnd! A dn PJ=0.0002 m=1 $X=46040 $Y=110300 $D=8
D110 A vdd! dn PJ=0.0002 m=1 $X=48360 $Y=-95300 $D=8
D111 A vdd! dn PJ=0.0002 m=1 $X=48360 $Y=114700 $D=8
D112 gnd! A dn PJ=0.0002 m=1 $X=50680 $Y=-99700 $D=8
D113 gnd! A dn PJ=0.0002 m=1 $X=50680 $Y=110300 $D=8
D114 A vdd! dn PJ=0.0002 m=1 $X=53000 $Y=-95300 $D=8
D115 A vdd! dn PJ=0.0002 m=1 $X=53000 $Y=114700 $D=8
D116 gnd! A dn PJ=0.0001 m=1 $X=55320 $Y=-99700 $D=8
D117 gnd! A dn PJ=0.0001 m=1 $X=55320 $Y=110300 $D=8
D118 A vdd! dn PJ=0.0001 m=1 $X=58500 $Y=4700 $D=8
D119 A vdd! dn PJ=0.0001 m=1 $X=58500 $Y=214700 $D=8
D120 gnd! A dn PJ=0.0002 m=1 $X=60820 $Y=-99700 $D=8
D121 gnd! A dn PJ=0.0002 m=1 $X=60820 $Y=110300 $D=8
D122 A vdd! dn PJ=0.0002 m=1 $X=63140 $Y=-95300 $D=8
D123 A vdd! dn PJ=0.0002 m=1 $X=63140 $Y=114700 $D=8
D124 gnd! A dn PJ=0.0002 m=1 $X=65460 $Y=-99700 $D=8
D125 gnd! A dn PJ=0.0002 m=1 $X=65460 $Y=110300 $D=8
D126 A vdd! dn PJ=0.0002 m=1 $X=67780 $Y=-95300 $D=8
D127 A vdd! dn PJ=0.0002 m=1 $X=67780 $Y=114700 $D=8
D128 gnd! A dn PJ=0.0001 m=1 $X=70100 $Y=-99700 $D=8
D129 gnd! A dn PJ=0.0001 m=1 $X=70100 $Y=110300 $D=8
D130 A vdd! dn PJ=0.0001 m=1 $X=73280 $Y=4700 $D=8
D131 A vdd! dn PJ=0.0001 m=1 $X=73280 $Y=214700 $D=8
D132 gnd! A dn PJ=0.0002 m=1 $X=75600 $Y=-99700 $D=8
D133 gnd! A dn PJ=0.0002 m=1 $X=75600 $Y=110300 $D=8
D134 A vdd! dn PJ=0.0002 m=1 $X=77920 $Y=-95300 $D=8
D135 A vdd! dn PJ=0.0002 m=1 $X=77920 $Y=114700 $D=8
D136 gnd! A dn PJ=0.0002 m=1 $X=80240 $Y=-99700 $D=8
D137 gnd! A dn PJ=0.0002 m=1 $X=80240 $Y=110300 $D=8
D138 A vdd! dn PJ=0.0002 m=1 $X=82560 $Y=-95300 $D=8
D139 A vdd! dn PJ=0.0002 m=1 $X=82560 $Y=114700 $D=8
D140 gnd! A dn PJ=0.0001 m=1 $X=84880 $Y=-99700 $D=8
D141 gnd! A dn PJ=0.0001 m=1 $X=84880 $Y=110300 $D=8
D142 A vdd! dn PJ=0.0001 m=1 $X=88060 $Y=4700 $D=8
D143 A vdd! dn PJ=0.0001 m=1 $X=88060 $Y=214700 $D=8
D144 gnd! A dn PJ=0.0002 m=1 $X=90380 $Y=-99700 $D=8
D145 gnd! A dn PJ=0.0002 m=1 $X=90380 $Y=110300 $D=8
D146 A vdd! dn PJ=0.0002 m=1 $X=92700 $Y=-95300 $D=8
D147 A vdd! dn PJ=0.0002 m=1 $X=92700 $Y=114700 $D=8
D148 gnd! A dn PJ=0.0002 m=1 $X=95020 $Y=-99700 $D=8
D149 gnd! A dn PJ=0.0002 m=1 $X=95020 $Y=110300 $D=8
D150 gnd! 30 dn PJ=5e-06 m=1 $X=1560 $Y=328560 $D=10
D151 30 vdd! dn PJ=5e-06 m=1 $X=1560 $Y=334960 $D=10
D152 gnd! 30 dn PJ=5e-06 m=1 $X=1560 $Y=329900 $D=11
D153 30 vdd! dn PJ=5e-06 m=1 $X=1560 $Y=332220 $D=11
X205 A 30 PAD $T=0 1440 0 0 $X=-5000 $Y=-235000
X210 gnd! vdd! cpoly_p_CDNS_5887047866568 $T=60980 317780 0 0 $X=60980 $Y=317780
X211 gnd! vdd! cpoly_p_CDNS_5887047866568 $T=65860 317780 0 0 $X=65860 $Y=317780
X212 gnd! vdd! cpoly_p_CDNS_5887047866568 $T=65860 326780 0 0 $X=65860 $Y=326780
X213 gnd! vdd! cpoly_p_CDNS_5887047866568 $T=70620 317780 0 0 $X=70620 $Y=317780
X214 gnd! vdd! cpoly_p_CDNS_5887047866568 $T=75500 317780 0 0 $X=75500 $Y=317780
X215 gnd! vdd! cpoly_p_CDNS_5887047866568 $T=75500 326780 0 0 $X=75500 $Y=326780
X216 gnd! vdd! cpoly_p_CDNS_5887047866568 $T=80260 317780 0 0 $X=80260 $Y=317780
X217 gnd! vdd! cpoly_p_CDNS_5887047866568 $T=85140 317780 0 0 $X=85140 $Y=317780
X218 gnd! vdd! cpoly_p_CDNS_5887047866568 $T=85140 326780 0 0 $X=85140 $Y=326780
X219 gnd! vdd! cpoly_p_CDNS_5887047866568 $T=89900 317780 0 0 $X=89900 $Y=317780
X220 gnd! vdd! cpoly_p_CDNS_5887047866568 $T=94780 317780 0 0 $X=94780 $Y=317780
X221 gnd! vdd! cpoly_p_CDNS_5887047866568 $T=94780 326780 0 0 $X=94780 $Y=326780
X222 gnd! 25 nSelect2 nmos_a_CDNS_5887047866521 $T=21720 329840 0 180 $X=20280 $Y=328340
X223 gnd! 25 nSelect1 nmos_a_CDNS_5887047866521 $T=23160 329840 0 180 $X=21720 $Y=328340
X224 vdd! gnd! cpoly_n_CDNS_5887047866570 $T=15960 336500 0 0 $X=15960 $Y=336500
X225 gnd! vdd! cpoly_p_CDNS_5887047866569 $T=15960 317780 0 0 $X=15960 $Y=317780
X226 vdd! gnd! cpoly_n_CDNS_5887047866571 $T=6800 336500 1 180 $X=1040 $Y=336500
.ENDS
***************************************
.SUBCKT ICV_83 1 2
** N=5 EP=2 IP=8 FDC=7152
X0 1 2 ICV_39 $T=0 0 0 0 $X=-360 $Y=-320
X1 1 2 ICV_39 $T=880960 0 0 0 $X=880600 $Y=-320
.ENDS
***************************************
.SUBCKT RingPad_AND3 In2 In1 Out In3 5 6 gnd! vdd!
** N=9 EP=8 IP=12 FDC=17
M0 5 In3 gnd! gnd! nmos_a L=2.4e-07 W=2.4e-06 AD=9.1e-13 AS=9.6e-13 PD=1.75e-06 PS=1.75e-06 w_cont=1.1e-06 nfing=1 source_num=2 $X=1180 $Y=13160 $D=1
M1 6 In2 5 5 nmos_a L=2.4e-07 W=2.4e-06 AD=1.4e-12 AS=6.24e-13 PD=3.5e-06 PS=1.75e-06 w_cont=1.1e-06 nfing=1 source_num=2 $X=2620 $Y=13160 $D=1
M2 9 In1 6 6 nmos_a L=2.4e-07 W=2.4e-06 AD=1.4e-12 AS=6.24e-13 PD=3.5e-06 PS=1.75e-06 w_cont=1.1e-06 nfing=1 source_num=2 $X=4820 $Y=13160 $D=1
M3 Out 9 gnd! gnd! nmos_a L=2.4e-07 W=4.8e-06 AD=1.0764e-12 AS=1.92e-12 PD=2.07e-06 PS=2.07e-06 w_cont=2.1e-06 nfing=1 source_num=2 $X=7580 $Y=9360 $D=1
M4 Out 9 gnd! gnd! nmos_a L=2.4e-07 W=4.8e-06 AD=1.0764e-12 AS=1.92e-12 PD=2.07e-06 PS=2.07e-06 w_cont=2.1e-06 nfing=1 source_num=2 $X=8340 $Y=9360 $D=1
M5 5 In3 gnd! gnd! nmos_a L=2.4e-07 W=2.4e-06 AD=9.1e-13 AS=9.6e-13 PD=1.75e-06 PS=1.75e-06 w_cont=1.1e-06 nfing=1 source_num=2 $X=420 $Y=13160 $D=1
M6 6 In2 5 5 nmos_a L=2.4e-07 W=2.4e-06 AD=1.4e-12 AS=6.24e-13 PD=3.5e-06 PS=1.75e-06 w_cont=1.1e-06 nfing=1 source_num=2 $X=3380 $Y=13160 $D=1
M7 9 In1 6 6 nmos_a L=2.4e-07 W=2.4e-06 AD=1.4e-12 AS=6.24e-13 PD=3.5e-06 PS=1.75e-06 w_cont=1.1e-06 nfing=1 source_num=2 $X=5580 $Y=13160 $D=1
M8 9 In3 vdd! vdd! pmos_a L=2.4e-07 W=2e-06 AD=6.76e-13 AS=1.3e-13 PD=1.3e-06 PS=1.3e-06 w_cont=6e-07 nfing=1 mmm=1 $X=1180 $Y=9360 $D=5
M9 9 In2 vdd! vdd! pmos_a L=2.4e-07 W=2e-06 AD=1.04e-12 AS=1.66e-13 PD=2.6e-06 PS=1.3e-06 w_cont=6e-07 nfing=1 mmm=1 $X=2620 $Y=9360 $D=5
M10 9 In2 vdd! vdd! pmos_a L=2.4e-07 W=2e-06 AD=1.04e-12 AS=1.66e-13 PD=2.6e-06 PS=1.3e-06 w_cont=6e-07 nfing=1 mmm=1 $X=3380 $Y=9360 $D=5
M11 9 In1 vdd! vdd! pmos_a L=2.4e-07 W=2e-06 AD=1.04e-12 AS=1.66e-13 PD=2.6e-06 PS=1.3e-06 w_cont=6e-07 nfing=1 mmm=1 $X=4820 $Y=9360 $D=5
M12 9 In1 vdd! vdd! pmos_a L=2.4e-07 W=2e-06 AD=1.04e-12 AS=1.66e-13 PD=2.6e-06 PS=1.3e-06 w_cont=6e-07 nfing=1 mmm=1 $X=5580 $Y=9360 $D=5
M13 Out 9 vdd! vdd! pmos_a L=2.4e-07 W=5.8e-06 AD=2.74097e-12 AS=3.12828e-13 PD=6.85241e-06 PS=3.42621e-06 w_cont=1.1e-06 nfing=1 mmm=1 $X=9780 $Y=9360 $D=5
M14 Out 9 vdd! vdd! pmos_a L=2.4e-07 W=5.8e-06 AD=1.78163e-12 AS=3.12828e-13 PD=3.42621e-06 PS=3.42621e-06 w_cont=1.1e-06 nfing=1 mmm=1 $X=10540 $Y=9360 $D=5
M15 Out 9 vdd! vdd! pmos_a L=2.4e-07 W=5.8e-06 AD=1.78163e-12 AS=2.47283e-13 PD=3.42621e-06 PS=3.42621e-06 w_cont=1.1e-06 nfing=1 mmm=1 $X=11300 $Y=9360 $D=5
M16 9 In3 vdd! vdd! pmos_a L=2.4e-07 W=2e-06 AD=6.76e-13 AS=1.3e-13 PD=1.3e-06 PS=1.3e-06 w_cont=6e-07 nfing=1 mmm=1 $X=420 $Y=9360 $D=5
.ENDS
***************************************
.SUBCKT PADIN_Adress nClk gnd! vdd! A nATD Adr
** N=24 EP=6 IP=164 FDC=120
M0 nATD 17 gnd! gnd! nmos_a L=2.4e-07 W=3.6e-06 AD=1.664e-12 AS=1.44e-12 PD=4.16e-06 PS=2.08e-06 w_cont=1.6e-06 nfing=1 source_num=2 $X=15140 $Y=324580 $D=1
M1 Adr 13 gnd! gnd! nmos_a L=2.4e-07 W=7.2e-06 AD=1.648e-12 AS=2.88e-12 PD=4.12e-06 PS=2.06e-06 w_cont=3.1e-06 nfing=1 source_num=2 $X=60100 $Y=319220 $D=1
M2 Adr 13 gnd! gnd! nmos_a L=2.4e-07 W=7.2e-06 AD=1.648e-12 AS=2.88e-12 PD=4.12e-06 PS=2.06e-06 w_cont=3.1e-06 nfing=1 source_num=2 $X=64840 $Y=319220 $D=1
M3 Adr 13 gnd! gnd! nmos_a L=2.4e-07 W=7.2e-06 AD=1.648e-12 AS=2.88e-12 PD=4.12e-06 PS=2.06e-06 w_cont=3.1e-06 nfing=1 source_num=2 $X=69740 $Y=319220 $D=1
M4 Adr 13 gnd! gnd! nmos_a L=2.4e-07 W=7.2e-06 AD=1.648e-12 AS=2.88e-12 PD=4.12e-06 PS=2.06e-06 w_cont=3.1e-06 nfing=1 source_num=2 $X=74480 $Y=319220 $D=1
M5 Adr 13 gnd! gnd! nmos_a L=2.4e-07 W=7.2e-06 AD=1.648e-12 AS=2.88e-12 PD=4.12e-06 PS=2.06e-06 w_cont=3.1e-06 nfing=1 source_num=2 $X=79380 $Y=319220 $D=1
M6 Adr 13 gnd! gnd! nmos_a L=2.4e-07 W=7.2e-06 AD=1.648e-12 AS=2.88e-12 PD=4.12e-06 PS=2.06e-06 w_cont=3.1e-06 nfing=1 source_num=2 $X=84120 $Y=319220 $D=1
M7 Adr 13 gnd! gnd! nmos_a L=2.4e-07 W=7.2e-06 AD=1.648e-12 AS=2.88e-12 PD=4.12e-06 PS=2.06e-06 w_cont=3.1e-06 nfing=1 source_num=2 $X=89020 $Y=319220 $D=1
M8 Adr 13 gnd! gnd! nmos_a L=2.4e-07 W=7.2e-06 AD=1.648e-12 AS=2.88e-12 PD=4.12e-06 PS=2.06e-06 w_cont=3.1e-06 nfing=1 source_num=2 $X=93760 $Y=319220 $D=1
M9 20 8 gnd! gnd! nmos_a L=2.4e-07 W=2.4e-06 AD=1.4e-12 AS=9.6e-13 PD=3.5e-06 PS=1.75e-06 w_cont=1.1e-06 nfing=1 source_num=2 $X=33840 $Y=326820 $D=1
M10 12 10 20 20 nmos_a L=2.4e-07 W=2.4e-06 AD=1.4e-12 AS=9.6e-13 PD=3.5e-06 PS=1.75e-06 w_cont=1.1e-06 nfing=1 source_num=2 $X=35280 $Y=326540 $D=1
M11 8 24 gnd! gnd! nmos_a L=2.4e-07 W=1.2e-06 AD=7.2e-13 AS=4.8e-13 PD=1.8e-06 PS=9e-07 w_cont=6e-07 nfing=1 source_num=2 $X=9380 $Y=325780 $D=1
M12 15 9 gnd! gnd! nmos_a L=2.4e-07 W=1.2e-06 AD=7.2e-13 AS=4.8e-13 PD=1.8e-06 PS=9e-07 w_cont=6e-07 nfing=1 source_num=2 $X=10820 $Y=325780 $D=1
M13 17 8 15 15 nmos_a L=2.4e-07 W=1.2e-06 AD=4.68e-13 AS=4.8e-13 PD=9e-07 PS=9e-07 w_cont=6e-07 nfing=1 source_num=2 $X=12320 $Y=328520 $D=1
M14 17 7 19 19 nmos_a L=2.4e-07 W=1.2e-06 AD=4.68e-13 AS=4.8e-13 PD=9e-07 PS=9e-07 w_cont=6e-07 nfing=1 source_num=2 $X=13080 $Y=328520 $D=1
M15 19 12 gnd! gnd! nmos_a L=2.4e-07 W=1.2e-06 AD=7.2e-13 AS=4.8e-13 PD=1.8e-06 PS=9e-07 w_cont=6e-07 nfing=1 source_num=2 $X=13700 $Y=325780 $D=1
M16 9 12 gnd! gnd! nmos_a L=2.4e-07 W=1.2e-06 AD=7.2e-13 AS=6.24e-13 PD=1.8e-06 PS=9e-07 w_cont=6e-07 nfing=1 source_num=2 $X=36680 $Y=327740 $D=1
M17 22 9 gnd! gnd! nmos_a L=2.4e-07 W=1.2e-06 AD=7.2e-13 AS=6.24e-13 PD=1.8e-06 PS=9e-07 w_cont=6e-07 nfing=1 source_num=2 $X=37440 $Y=327740 $D=1
M18 12 11 22 22 nmos_a L=2.4e-07 W=1.2e-06 AD=7.2e-13 AS=4.8e-13 PD=1.8e-06 PS=9e-07 w_cont=6e-07 nfing=1 source_num=2 $X=38880 $Y=327420 $D=1
M19 10 11 gnd! gnd! nmos_a L=2.4e-07 W=1.2e-06 AD=7.2e-13 AS=4.8e-13 PD=1.8e-06 PS=9e-07 w_cont=6e-07 nfing=1 source_num=2 $X=40280 $Y=327420 $D=1
M20 11 nClk gnd! gnd! nmos_a L=2.4e-07 W=1.2e-06 AD=7.2e-13 AS=4.8e-13 PD=1.8e-06 PS=9e-07 w_cont=6e-07 nfing=1 source_num=2 $X=41720 $Y=327420 $D=1
M21 7 8 gnd! gnd! nmos_a L=2.4e-07 W=4.8e-07 AD=4.32e-13 AS=1.92e-13 PD=1.08e-06 PS=5.4e-07 w_cont=6e-07 nfing=1 source_num=2 $X=12260 $Y=325980 $D=1
M22 13 12 gnd! gnd! nmos_a L=2.4e-07 W=3.6e-06 AD=1.664e-12 AS=1.44e-12 PD=4.16e-06 PS=2.08e-06 w_cont=1.6e-06 nfing=1 source_num=2 $X=47800 $Y=327560 $D=1
M23 13 12 gnd! gnd! nmos_a L=2.4e-07 W=3.6e-06 AD=1.664e-12 AS=1.44e-12 PD=4.16e-06 PS=2.08e-06 w_cont=1.6e-06 nfing=1 source_num=2 $X=53880 $Y=327560 $D=1
M24 18 9 vdd! vdd! pmos_a L=2.4e-07 W=2e-06 AD=1.04e-12 AS=1.3e-13 PD=2.6e-06 PS=1.3e-06 w_cont=6e-07 nfing=1 mmm=1 $X=13640 $Y=334500 $D=5
M25 nATD 17 vdd! vdd! pmos_a L=2.4e-07 W=5.76e-06 AD=2.744e-12 AS=2.488e-13 PD=6.86e-06 PS=3.43e-06 w_cont=1.1e-06 nfing=1 mmm=1 $X=15140 $Y=330600 $D=5
M26 Adr 13 vdd! vdd! pmos_a L=2.4e-07 W=1.1e-05 AD=2.63913e-12 AS=1.96364e-13 PD=6.59782e-06 PS=3.29891e-06 w_cont=1.6e-06 nfing=1 mmm=1 $X=60100 $Y=330700 $D=5
M27 Adr 13 vdd! vdd! pmos_a L=2.4e-07 W=1.1e-05 AD=2.63913e-12 AS=1.96364e-13 PD=6.59782e-06 PS=3.29891e-06 w_cont=1.6e-06 nfing=1 mmm=1 $X=64840 $Y=330700 $D=5
M28 Adr 13 vdd! vdd! pmos_a L=2.4e-07 W=1.1e-05 AD=2.63913e-12 AS=1.96364e-13 PD=6.59782e-06 PS=3.29891e-06 w_cont=1.6e-06 nfing=1 mmm=1 $X=69740 $Y=330700 $D=5
M29 Adr 13 vdd! vdd! pmos_a L=2.4e-07 W=1.088e-05 AD=2.64282e-12 AS=1.98212e-13 PD=6.60706e-06 PS=3.30353e-06 w_cont=1.6e-06 nfing=1 mmm=1 $X=74480 $Y=330820 $D=5
M30 Adr 13 vdd! vdd! pmos_a L=2.4e-07 W=1.1e-05 AD=2.63913e-12 AS=1.96364e-13 PD=6.59782e-06 PS=3.29891e-06 w_cont=1.6e-06 nfing=1 mmm=1 $X=79380 $Y=330700 $D=5
M31 Adr 13 vdd! vdd! pmos_a L=2.4e-07 W=1.1e-05 AD=2.63913e-12 AS=1.96364e-13 PD=6.59782e-06 PS=3.29891e-06 w_cont=1.6e-06 nfing=1 mmm=1 $X=84120 $Y=330700 $D=5
M32 Adr 13 vdd! vdd! pmos_a L=2.4e-07 W=1.1e-05 AD=2.63913e-12 AS=1.96364e-13 PD=6.59782e-06 PS=3.29891e-06 w_cont=1.6e-06 nfing=1 mmm=1 $X=89020 $Y=330700 $D=5
M33 Adr 13 vdd! vdd! pmos_a L=2.4e-07 W=1.1e-05 AD=2.63913e-12 AS=1.96364e-13 PD=6.59782e-06 PS=3.29891e-06 w_cont=1.6e-06 nfing=1 mmm=1 $X=93760 $Y=330700 $D=5
M34 13 12 vdd! vdd! pmos_a L=2.4e-07 W=5.76e-06 AD=2.744e-12 AS=2.488e-13 PD=6.86e-06 PS=3.43e-06 w_cont=1.1e-06 nfing=1 mmm=1 $X=46400 $Y=327560 $D=5
M35 13 12 vdd! vdd! pmos_a L=2.4e-07 W=5.76e-06 AD=2.744e-12 AS=2.488e-13 PD=6.86e-06 PS=3.43e-06 w_cont=1.1e-06 nfing=1 mmm=1 $X=52480 $Y=327560 $D=5
M36 14 14 vdd! vdd! pmos_a L=2.4e-07 W=2e-06 AD=6.76e-13 AS=1.3e-13 PD=1.3e-06 PS=1.3e-06 w_cont=6e-07 nfing=1 mmm=1 $X=9240 $Y=334300 $D=5
M37 14 14 vdd! vdd! pmos_a L=2.4e-07 W=2e-06 AD=6.76e-13 AS=1.66e-13 PD=1.3e-06 PS=1.3e-06 w_cont=6e-07 nfing=1 mmm=1 $X=10000 $Y=334300 $D=5
M38 16 12 vdd! vdd! pmos_a L=2.4e-07 W=2e-06 AD=1.04e-12 AS=1.66e-13 PD=2.6e-06 PS=1.3e-06 w_cont=6e-07 nfing=1 mmm=1 $X=10760 $Y=334300 $D=5
M39 17 8 16 16 pmos_a L=2.4e-07 W=2e-06 AD=6.76e-13 AS=1.3e-13 PD=1.3e-06 PS=1.3e-06 w_cont=6e-07 nfing=1 mmm=1 $X=12320 $Y=331000 $D=5
M40 17 7 18 18 pmos_a L=2.4e-07 W=2e-06 AD=6.76e-13 AS=1.3e-13 PD=1.3e-06 PS=1.3e-06 w_cont=6e-07 nfing=1 mmm=1 $X=13080 $Y=331000 $D=5
M41 9 12 vdd! vdd! pmos_a L=2.4e-07 W=2e-06 AD=1.04e-12 AS=1.66e-13 PD=2.6e-06 PS=1.3e-06 w_cont=6e-07 nfing=1 mmm=1 $X=36680 $Y=330700 $D=5
M42 23 9 vdd! vdd! pmos_a L=2.4e-07 W=2e-06 AD=1.04e-12 AS=1.66e-13 PD=2.6e-06 PS=1.3e-06 w_cont=6e-07 nfing=1 mmm=1 $X=37440 $Y=330700 $D=5
M43 12 10 23 23 pmos_a L=2.4e-07 W=2e-06 AD=1.04e-12 AS=1.3e-13 PD=2.6e-06 PS=1.3e-06 w_cont=6e-07 nfing=1 mmm=1 $X=38880 $Y=330200 $D=5
M44 10 11 vdd! vdd! pmos_a L=2.4e-07 W=2e-06 AD=1.04e-12 AS=1.3e-13 PD=2.6e-06 PS=1.3e-06 w_cont=6e-07 nfing=1 mmm=1 $X=40280 $Y=330200 $D=5
M45 11 nClk vdd! vdd! pmos_a L=2.4e-07 W=2e-06 AD=1.04e-12 AS=1.3e-13 PD=2.6e-06 PS=1.3e-06 w_cont=6e-07 nfing=1 mmm=1 $X=41720 $Y=331700 $D=5
M46 7 8 vdd! vdd! pmos_a L=2.4e-07 W=1e-06 AD=6.4e-13 AS=1.25e-13 PD=1.6e-06 PS=8e-07 w_cont=6e-07 nfing=1 mmm=1 $X=12200 $Y=335000 $D=5
M47 14 7 vdd! vdd! pmos_a L=2.4e-07 W=4e-06 AD=1.84e-12 AS=1.4e-13 PD=4.6e-06 PS=2.3e-06 w_cont=6e-07 nfing=1 mmm=1 $X=8800 $Y=329000 $D=5
M48 8 24 14 14 pmos_a L=2.4e-07 W=4e-06 AD=1.84e-12 AS=1.4e-13 PD=4.6e-06 PS=2.3e-06 w_cont=6e-07 nfing=1 mmm=1 $X=10240 $Y=328320 $D=5
M49 21 8 vdd! vdd! pmos_a L=2.4e-07 W=4e-06 AD=1.84e-12 AS=1.4e-13 PD=4.6e-06 PS=2.3e-06 w_cont=6e-07 nfing=1 mmm=1 $X=33840 $Y=331020 $D=5
M50 12 11 21 21 pmos_a L=2.4e-07 W=4e-06 AD=1.84e-12 AS=1.4e-13 PD=4.6e-06 PS=2.3e-06 w_cont=6e-07 nfing=1 mmm=1 $X=35280 $Y=331020 $D=5
M51 vdd! gnd! vdd! cpoly_n w=6e-06 l=2e-06 c=7.5402e-14 as=2.4e-13 ad=2.304e-12 ps=2.88e-06 pd=4.86761e-06 sim_w=5.76e-06 m_per_maxw=1.04167 numb_sub_cont=3 nfing=1 $X=30600 $Y=328520 $D=22
M52 vdd! gnd! vdd! cpoly_n w=6e-06 l=2e-06 c=7.5402e-14 as=2.4e-13 ad=2.304e-12 ps=2.88e-06 pd=4.86761e-06 sim_w=5.76e-06 m_per_maxw=1.04167 numb_sub_cont=3 nfing=1 $X=43200 $Y=328200 $D=22
M53 vdd! gnd! vdd! cpoly_n w=6e-06 l=2e-06 c=7.5402e-14 as=2.4e-13 ad=2.304e-12 ps=2.88e-06 pd=4.86761e-06 sim_w=5.76e-06 m_per_maxw=1.04167 numb_sub_cont=3 nfing=1 $X=49280 $Y=328200 $D=22
M54 vdd! gnd! vdd! cpoly_n w=6e-06 l=2e-06 c=7.5402e-14 as=2.4e-13 ad=2.304e-12 ps=2.88e-06 pd=4.86761e-06 sim_w=5.76e-06 m_per_maxw=1.04167 numb_sub_cont=3 nfing=1 $X=55360 $Y=328200 $D=22
M55 vdd! gnd! vdd! cpoly_n w=6e-06 l=2e-06 c=7.5402e-14 as=2.4e-13 ad=2.304e-12 ps=2.88e-06 pd=4.86761e-06 sim_w=5.76e-06 m_per_maxw=1.04167 numb_sub_cont=3 nfing=1 $X=61600 $Y=328200 $D=22
M56 vdd! gnd! vdd! cpoly_n w=6e-06 l=2e-06 c=7.5402e-14 as=2.4e-13 ad=2.304e-12 ps=2.88e-06 pd=4.86761e-06 sim_w=5.76e-06 m_per_maxw=1.04167 numb_sub_cont=3 nfing=1 $X=61600 $Y=336700 $D=22
M57 vdd! gnd! vdd! cpoly_n w=6e-06 l=2e-06 c=7.5402e-14 as=2.4e-13 ad=2.304e-12 ps=2.88e-06 pd=4.86761e-06 sim_w=5.76e-06 m_per_maxw=1.04167 numb_sub_cont=3 nfing=1 $X=66480 $Y=336700 $D=22
M58 vdd! gnd! vdd! cpoly_n w=6e-06 l=2e-06 c=7.5402e-14 as=2.4e-13 ad=2.304e-12 ps=2.88e-06 pd=4.86761e-06 sim_w=5.76e-06 m_per_maxw=1.04167 numb_sub_cont=3 nfing=1 $X=71240 $Y=328200 $D=22
M59 vdd! gnd! vdd! cpoly_n w=6e-06 l=2e-06 c=7.5402e-14 as=2.4e-13 ad=2.304e-12 ps=2.88e-06 pd=4.86761e-06 sim_w=5.76e-06 m_per_maxw=1.04167 numb_sub_cont=3 nfing=1 $X=71240 $Y=336700 $D=22
M60 vdd! gnd! vdd! cpoly_n w=6e-06 l=2e-06 c=7.5402e-14 as=2.4e-13 ad=2.304e-12 ps=2.88e-06 pd=4.86761e-06 sim_w=5.76e-06 m_per_maxw=1.04167 numb_sub_cont=3 nfing=1 $X=76120 $Y=336700 $D=22
M61 vdd! gnd! vdd! cpoly_n w=6e-06 l=2e-06 c=7.5402e-14 as=2.4e-13 ad=2.304e-12 ps=2.88e-06 pd=4.86761e-06 sim_w=5.76e-06 m_per_maxw=1.04167 numb_sub_cont=3 nfing=1 $X=80880 $Y=328200 $D=22
M62 vdd! gnd! vdd! cpoly_n w=6e-06 l=2e-06 c=7.5402e-14 as=2.4e-13 ad=2.304e-12 ps=2.88e-06 pd=4.86761e-06 sim_w=5.76e-06 m_per_maxw=1.04167 numb_sub_cont=3 nfing=1 $X=80880 $Y=336700 $D=22
M63 vdd! gnd! vdd! cpoly_n w=6e-06 l=2e-06 c=7.5402e-14 as=2.4e-13 ad=2.304e-12 ps=2.88e-06 pd=4.86761e-06 sim_w=5.76e-06 m_per_maxw=1.04167 numb_sub_cont=3 nfing=1 $X=85760 $Y=336700 $D=22
M64 vdd! gnd! vdd! cpoly_n w=6e-06 l=2e-06 c=7.5402e-14 as=2.4e-13 ad=2.304e-12 ps=2.88e-06 pd=4.86761e-06 sim_w=5.76e-06 m_per_maxw=1.04167 numb_sub_cont=3 nfing=1 $X=90520 $Y=328200 $D=22
M65 vdd! gnd! vdd! cpoly_n w=6e-06 l=2e-06 c=7.5402e-14 as=2.4e-13 ad=2.304e-12 ps=2.88e-06 pd=4.86761e-06 sim_w=5.76e-06 m_per_maxw=1.04167 numb_sub_cont=3 nfing=1 $X=90520 $Y=336700 $D=22
M66 vdd! gnd! vdd! cpoly_n w=6e-06 l=2e-06 c=7.5402e-14 as=2.4e-13 ad=2.304e-12 ps=2.88e-06 pd=4.86761e-06 sim_w=5.76e-06 m_per_maxw=1.04167 numb_sub_cont=3 nfing=1 $X=95400 $Y=336700 $D=22
D67 gnd! 24 dn PJ=5e-06 m=1 $X=1560 $Y=328560 $D=10
D68 24 vdd! dn PJ=5e-06 m=1 $X=1560 $Y=334960 $D=10
D69 gnd! 24 dn PJ=5e-06 m=1 $X=1560 $Y=329900 $D=11
D70 24 vdd! dn PJ=5e-06 m=1 $X=1560 $Y=332220 $D=11
X115 A 24 PAD $T=0 1440 0 0 $X=-5000 $Y=-235000
X120 gnd! vdd! cpoly_p_CDNS_5887047866568 $T=60980 317780 0 0 $X=60980 $Y=317780
X121 gnd! vdd! cpoly_p_CDNS_5887047866568 $T=65860 317780 0 0 $X=65860 $Y=317780
X122 gnd! vdd! cpoly_p_CDNS_5887047866568 $T=65860 326780 0 0 $X=65860 $Y=326780
X123 gnd! vdd! cpoly_p_CDNS_5887047866568 $T=70620 317780 0 0 $X=70620 $Y=317780
X124 gnd! vdd! cpoly_p_CDNS_5887047866568 $T=75500 317780 0 0 $X=75500 $Y=317780
X125 gnd! vdd! cpoly_p_CDNS_5887047866568 $T=75500 326780 0 0 $X=75500 $Y=326780
X126 gnd! vdd! cpoly_p_CDNS_5887047866568 $T=80260 317780 0 0 $X=80260 $Y=317780
X127 gnd! vdd! cpoly_p_CDNS_5887047866568 $T=85140 317780 0 0 $X=85140 $Y=317780
X128 gnd! vdd! cpoly_p_CDNS_5887047866568 $T=85140 326780 0 0 $X=85140 $Y=326780
X129 gnd! vdd! cpoly_p_CDNS_5887047866568 $T=89900 317780 0 0 $X=89900 $Y=317780
X130 gnd! vdd! cpoly_p_CDNS_5887047866568 $T=94780 317780 0 0 $X=94780 $Y=317780
X131 gnd! vdd! cpoly_p_CDNS_5887047866568 $T=94780 326780 0 0 $X=94780 $Y=326780
X132 vdd! gnd! cpoly_n_CDNS_5887047866570 $T=15960 336500 0 0 $X=15960 $Y=336500
X133 gnd! vdd! cpoly_p_CDNS_5887047866569 $T=15960 317780 0 0 $X=15960 $Y=317780
X134 vdd! gnd! cpoly_n_CDNS_5887047866571 $T=6800 336500 1 180 $X=1040 $Y=336500
.ENDS
***************************************
.SUBCKT ICV_84 1 2 3
** N=3 EP=3 IP=4 FDC=2
D0 2 1 dn PJ=0.00041 m=1 $X=-460 $Y=0 $D=9
D1 3 2 dn PJ=0.00041 m=1 $X=2040 $Y=0 $D=9
.ENDS
***************************************
.SUBCKT ICV_85 1 2 3
** N=3 EP=3 IP=6 FDC=4
X0 1 2 3 ICV_31 $T=5000 0 0 0 $X=4360 $Y=-300
X1 3 2 1 ICV_84 $T=0 0 0 0 $X=-640 $Y=-300
.ENDS
***************************************
.SUBCKT ICV_86 1 2 3
** N=3 EP=3 IP=6 FDC=8
X0 3 2 1 ICV_85 $T=0 0 0 0 $X=-640 $Y=-300
X1 3 2 1 ICV_85 $T=10000 0 0 0 $X=9360 $Y=-300
.ENDS
***************************************
.SUBCKT GND_PAD GND_PAD VDD_PAD gnd! vdd!
** N=8 EP=4 IP=21 FDC=115
D0 GND_PAD VDD_PAD dn PJ=0.00041 m=1 $X=94260 $Y=-99700 $D=9
X1 vdd! gnd! cpoly_n_CDNS_588704786651 $T=520 333340 0 0 $X=520 $Y=333340
X2 gnd! vdd! cpoly_p_CDNS_588704786650 $T=520 320500 0 0 $X=520 $Y=320500
X4 gnd! GND_PAD VDD_PAD ICV_85 $T=84720 -99700 0 0 $X=84080 $Y=-100000
X5 VDD_PAD GND_PAD gnd! ICV_86 $T=4720 -99700 0 0 $X=4080 $Y=-100000
X6 VDD_PAD GND_PAD gnd! ICV_86 $T=24720 -99700 0 0 $X=24080 $Y=-100000
X7 VDD_PAD GND_PAD gnd! ICV_86 $T=44720 -99700 0 0 $X=44080 $Y=-100000
X8 VDD_PAD GND_PAD gnd! ICV_86 $T=64720 -99700 0 0 $X=64080 $Y=-100000
.ENDS
***************************************
.SUBCKT nOE_16 Bit_16 Bit_32 gnd! nOE Out vdd!
** N=10 EP=6 IP=0 FDC=10
M0 Out 8 gnd! gnd! nmos_a L=2.4e-07 W=4.8e-07 AD=4.32e-13 AS=1.92e-13 PD=1.08e-06 PS=5.4e-07 w_cont=6e-07 nfing=1 source_num=2 $X=1040 $Y=640 $D=1
M1 8 nOE gnd! gnd! nmos_a L=2.4e-07 W=4.8e-07 AD=4.32e-13 AS=1.92e-13 PD=1.08e-06 PS=5.4e-07 w_cont=6e-07 nfing=1 source_num=2 $X=2480 $Y=640 $D=1
M2 8 10 gnd! gnd! nmos_a L=2.4e-07 W=4.8e-07 AD=4.32e-13 AS=1.92e-13 PD=1.08e-06 PS=5.4e-07 w_cont=6e-07 nfing=1 source_num=2 $X=3920 $Y=640 $D=1
M3 10 Bit_16 gnd! gnd! nmos_a L=2.4e-07 W=4.8e-07 AD=4.32e-13 AS=1.92e-13 PD=1.08e-06 PS=5.4e-07 w_cont=6e-07 nfing=1 source_num=2 $X=5360 $Y=640 $D=1
M4 10 Bit_32 gnd! gnd! nmos_a L=2.4e-07 W=4.8e-07 AD=4.32e-13 AS=1.92e-13 PD=1.08e-06 PS=5.4e-07 w_cont=6e-07 nfing=1 source_num=2 $X=6800 $Y=640 $D=1
M5 Out 8 vdd! vdd! pmos_a L=2.4e-07 W=1e-06 AD=6.4e-13 AS=1.25e-13 PD=1.6e-06 PS=8e-07 w_cont=6e-07 nfing=1 mmm=1 $X=1040 $Y=2960 $D=5
M6 7 nOE vdd! vdd! pmos_a L=2.4e-07 W=1e-06 AD=6.4e-13 AS=1.25e-13 PD=1.6e-06 PS=8e-07 w_cont=6e-07 nfing=1 mmm=1 $X=2480 $Y=2960 $D=5
M7 8 10 7 7 pmos_a L=2.4e-07 W=1e-06 AD=6.4e-13 AS=1.25e-13 PD=1.6e-06 PS=8e-07 w_cont=6e-07 nfing=1 mmm=1 $X=3920 $Y=2960 $D=5
M8 9 Bit_16 vdd! vdd! pmos_a L=2.4e-07 W=1e-06 AD=6.4e-13 AS=1.25e-13 PD=1.6e-06 PS=8e-07 w_cont=6e-07 nfing=1 mmm=1 $X=5360 $Y=2960 $D=5
M9 10 Bit_32 9 9 pmos_a L=2.4e-07 W=1e-06 AD=6.4e-13 AS=1.25e-13 PD=1.6e-06 PS=8e-07 w_cont=6e-07 nfing=1 mmm=1 $X=6800 $Y=2960 $D=5
.ENDS
***************************************
.SUBCKT cpoly_n_CDNS_5887047866566 1 2
** N=2 EP=2 IP=0 FDC=3
M0 1 2 1 cpoly_n w=6e-06 l=2e-06 c=7.5402e-14 as=2.4e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.4338e-06 sim_w=5.76e-06 m_per_maxw=1.04167 numb_sub_cont=3 nfing=1 $X=620 $Y=200 $D=22
M1 1 2 1 cpoly_n w=6e-06 l=2e-06 c=7.5402e-14 as=3.0336e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.4338e-06 sim_w=5.76e-06 m_per_maxw=1.04167 numb_sub_cont=3 nfing=1 $X=3140 $Y=200 $D=22
M2 1 2 1 cpoly_n w=6e-06 l=2e-06 c=7.5402e-14 as=3.0336e-13 ad=2.304e-12 ps=2.88e-06 pd=4.86761e-06 sim_w=5.76e-06 m_per_maxw=1.04167 numb_sub_cont=3 nfing=1 $X=5660 $Y=200 $D=22
.ENDS
***************************************
.SUBCKT pmos_a_CDNS_5887047866512
** N=3 EP=0 IP=0 FDC=0
*.SEEDPROM
.ENDS
***************************************
.SUBCKT ICV_87 1 2 3 4
** N=4 EP=4 IP=6 FDC=2
M0 2 4 1 1 nmos_a L=2.4e-07 W=2.4e-06 AD=1.4e-12 AS=9.6e-13 PD=3.5e-06 PS=1.75e-06 w_cont=1.1e-06 nfing=1 source_num=2 $X=620 $Y=200 $D=1
M1 2 4 3 3 pmos_a L=2.4e-07 W=4.5e-06 AD=2.04e-12 AS=1.425e-13 PD=5.1e-06 PS=2.55e-06 w_cont=6e-07 nfing=1 mmm=1 $X=620 $Y=4600 $D=5
.ENDS
***************************************
.SUBCKT PADIN_OE gnd! vdd! OEN WEN CE nOE nOE_Master
** N=17 EP=7 IP=88 FDC=212
M0 8 10 gnd! gnd! nmos_a L=2.4e-07 W=1.2e-06 AD=7.2e-13 AS=6.24e-13 PD=1.8e-06 PS=9e-07 w_cont=6e-07 nfing=1 source_num=2 $X=10960 $Y=328200 $D=1
M1 14 WEN 12 12 nmos_a L=2.4e-07 W=1e-06 AD=6.4e-13 AS=4e-13 PD=1.6e-06 PS=8e-07 w_cont=6e-07 nfing=1 source_num=2 $X=12640 $Y=328820 $D=1
M2 12 CE 13 13 nmos_a L=2.4e-07 W=1e-06 AD=6.4e-13 AS=4e-13 PD=1.6e-06 PS=8e-07 w_cont=6e-07 nfing=1 source_num=2 $X=14080 $Y=328820 $D=1
M3 13 16 gnd! gnd! nmos_a L=2.4e-07 W=1e-06 AD=6.4e-13 AS=5.2e-13 PD=1.6e-06 PS=8e-07 w_cont=6e-07 nfing=1 source_num=2 $X=15520 $Y=328820 $D=1
M4 15 14 gnd! gnd! nmos_a L=2.4e-07 W=1e-06 AD=6.4e-13 AS=5.2e-13 PD=1.6e-06 PS=8e-07 w_cont=6e-07 nfing=1 source_num=2 $X=16280 $Y=328820 $D=1
M5 16 nOE 15 15 nmos_a L=2.4e-07 W=1e-06 AD=6.4e-13 AS=4e-13 PD=1.6e-06 PS=8e-07 w_cont=6e-07 nfing=1 source_num=2 $X=17720 $Y=328820 $D=1
M6 10 14 gnd! gnd! nmos_a L=2.4e-07 W=1.2e-06 AD=7.2e-13 AS=6.24e-13 PD=1.8e-06 PS=9e-07 w_cont=6e-07 nfing=1 source_num=2 $X=10200 $Y=328200 $D=1
M7 10 17 gnd! gnd! nmos_a L=2.4e-07 W=4.8e-07 AD=4.32e-13 AS=1.92e-13 PD=1.08e-06 PS=5.4e-07 w_cont=6e-07 nfing=1 source_num=2 $X=8800 $Y=328200 $D=1
M8 11 8 vdd! vdd! pmos_a L=4e-07 W=4.8e-07 AD=4.32e-13 AS=1.224e-13 PD=1.08e-06 PS=5.4e-07 w_cont=6e-07 nfing=1 mmm=1 $X=10240 $Y=333300 $D=5
M9 8 10 vdd! vdd! pmos_a L=2.4e-07 W=2e-06 AD=1.04e-12 AS=1.3e-13 PD=2.6e-06 PS=1.3e-06 w_cont=6e-07 nfing=1 mmm=1 $X=11840 $Y=332300 $D=5
M10 14 WEN vdd! vdd! pmos_a L=2.4e-07 W=7e-07 AD=3.38e-13 AS=1.295e-13 PD=6.5e-07 PS=6.5e-07 w_cont=6e-07 nfing=1 mmm=1 $X=13320 $Y=331860 $D=5
M11 14 CE vdd! vdd! pmos_a L=2.4e-07 W=7e-07 AD=3.38e-13 AS=1.595e-13 PD=6.5e-07 PS=6.5e-07 w_cont=6e-07 nfing=1 mmm=1 $X=14080 $Y=331860 $D=5
M12 14 16 vdd! vdd! pmos_a L=2.4e-07 W=7e-07 AD=5.2e-13 AS=1.595e-13 PD=1.3e-06 PS=6.5e-07 w_cont=6e-07 nfing=1 mmm=1 $X=14840 $Y=331860 $D=5
M13 16 14 vdd! vdd! pmos_a L=2.4e-07 W=1e-06 AD=6.4e-13 AS=1.61e-13 PD=1.6e-06 PS=8e-07 w_cont=6e-07 nfing=1 mmm=1 $X=16960 $Y=332120 $D=5
M14 16 nOE vdd! vdd! pmos_a L=2.4e-07 W=1e-06 AD=6.4e-13 AS=1.61e-13 PD=1.6e-06 PS=8e-07 w_cont=6e-07 nfing=1 mmm=1 $X=17720 $Y=332120 $D=5
M15 10 17 11 11 pmos_a L=2.4e-07 W=1e-06 AD=6.4e-13 AS=1.25e-13 PD=1.6e-06 PS=8e-07 w_cont=6e-07 nfing=1 mmm=1 $X=8800 $Y=330180 $D=5
M16 11 14 vdd! vdd! pmos_a L=2.4e-07 W=1e-06 AD=6.4e-13 AS=1.25e-13 PD=1.6e-06 PS=8e-07 w_cont=6e-07 nfing=1 mmm=1 $X=8820 $Y=332980 $D=5
M17 vdd! gnd! vdd! cpoly_n w=6e-06 l=2e-06 c=7.5402e-14 as=2.4e-13 ad=2.304e-12 ps=2.88e-06 pd=4.86761e-06 sim_w=5.76e-06 m_per_maxw=1.04167 numb_sub_cont=3 nfing=1 $X=20680 $Y=328200 $D=22
M18 vdd! gnd! vdd! cpoly_n w=6e-06 l=2e-06 c=7.5402e-14 as=3.0336e-13 ad=2.304e-12 ps=2.88e-06 pd=4.86761e-06 sim_w=5.76e-06 m_per_maxw=1.04167 numb_sub_cont=3 nfing=1 $X=25280 $Y=328200 $D=22
M19 vdd! gnd! vdd! cpoly_n w=6e-06 l=2e-06 c=7.5402e-14 as=3.0336e-13 ad=2.304e-12 ps=2.88e-06 pd=4.86761e-06 sim_w=5.76e-06 m_per_maxw=1.04167 numb_sub_cont=3 nfing=1 $X=27800 $Y=328200 $D=22
M20 vdd! gnd! vdd! cpoly_n w=6e-06 l=2e-06 c=7.5402e-14 as=2.4e-13 ad=2.304e-12 ps=2.88e-06 pd=4.86761e-06 sim_w=5.76e-06 m_per_maxw=1.04167 numb_sub_cont=3 nfing=1 $X=32440 $Y=328200 $D=22
M21 vdd! gnd! vdd! cpoly_n w=6e-06 l=2e-06 c=7.5402e-14 as=2.4e-13 ad=2.304e-12 ps=2.88e-06 pd=4.86761e-06 sim_w=5.76e-06 m_per_maxw=1.04167 numb_sub_cont=3 nfing=1 $X=37080 $Y=328200 $D=22
M22 vdd! gnd! vdd! cpoly_n w=6e-06 l=2e-06 c=7.5402e-14 as=2.4e-13 ad=2.304e-12 ps=2.88e-06 pd=4.86761e-06 sim_w=5.76e-06 m_per_maxw=1.04167 numb_sub_cont=3 nfing=1 $X=41720 $Y=328200 $D=22
M23 vdd! gnd! vdd! cpoly_n w=6e-06 l=2e-06 c=7.5402e-14 as=2.4e-13 ad=2.304e-12 ps=2.88e-06 pd=4.86761e-06 sim_w=5.76e-06 m_per_maxw=1.04167 numb_sub_cont=3 nfing=1 $X=46360 $Y=328200 $D=22
M24 vdd! gnd! vdd! cpoly_n w=6e-06 l=2e-06 c=7.5402e-14 as=2.4e-13 ad=2.304e-12 ps=2.88e-06 pd=4.86761e-06 sim_w=5.76e-06 m_per_maxw=1.04167 numb_sub_cont=3 nfing=1 $X=51000 $Y=328200 $D=22
M25 vdd! gnd! vdd! cpoly_n w=6e-06 l=2e-06 c=7.5402e-14 as=2.4e-13 ad=2.304e-12 ps=2.88e-06 pd=4.86761e-06 sim_w=5.76e-06 m_per_maxw=1.04167 numb_sub_cont=3 nfing=1 $X=55640 $Y=328200 $D=22
M26 vdd! gnd! vdd! cpoly_n w=6e-06 l=2e-06 c=7.5402e-14 as=2.4e-13 ad=2.304e-12 ps=2.88e-06 pd=4.86761e-06 sim_w=5.76e-06 m_per_maxw=1.04167 numb_sub_cont=3 nfing=1 $X=60280 $Y=328200 $D=22
D27 OEN vdd! dn PJ=0.0002 m=1 $X=4020 $Y=-95300 $D=9
D28 OEN vdd! dn PJ=0.0002 m=1 $X=4020 $Y=114700 $D=9
D29 gnd! OEN dn PJ=0.0002 m=1 $X=6340 $Y=-99700 $D=9
D30 gnd! OEN dn PJ=0.0002 m=1 $X=6340 $Y=110300 $D=9
D31 OEN vdd! dn PJ=0.0002 m=1 $X=8660 $Y=-95300 $D=9
D32 OEN vdd! dn PJ=0.0002 m=1 $X=8660 $Y=114700 $D=9
D33 gnd! OEN dn PJ=0.0001 m=1 $X=10980 $Y=-99700 $D=9
D34 gnd! OEN dn PJ=0.0001 m=1 $X=10980 $Y=110300 $D=9
D35 OEN vdd! dn PJ=0.0001 m=1 $X=14160 $Y=4700 $D=9
D36 OEN vdd! dn PJ=0.0001 m=1 $X=14160 $Y=214700 $D=9
D37 gnd! OEN dn PJ=0.0002 m=1 $X=16480 $Y=-99700 $D=9
D38 gnd! OEN dn PJ=0.0002 m=1 $X=16480 $Y=110300 $D=9
D39 OEN vdd! dn PJ=0.0002 m=1 $X=18800 $Y=-95300 $D=9
D40 OEN vdd! dn PJ=0.0002 m=1 $X=18800 $Y=114700 $D=9
D41 gnd! OEN dn PJ=0.0002 m=1 $X=21120 $Y=-99700 $D=9
D42 gnd! OEN dn PJ=0.0002 m=1 $X=21120 $Y=110300 $D=9
D43 OEN vdd! dn PJ=0.0002 m=1 $X=23440 $Y=-95300 $D=9
D44 OEN vdd! dn PJ=0.0002 m=1 $X=23440 $Y=114700 $D=9
D45 gnd! OEN dn PJ=0.0001 m=1 $X=25760 $Y=-99700 $D=9
D46 gnd! OEN dn PJ=0.0001 m=1 $X=25760 $Y=110300 $D=9
D47 OEN vdd! dn PJ=0.0001 m=1 $X=28940 $Y=4700 $D=9
D48 OEN vdd! dn PJ=0.0001 m=1 $X=28940 $Y=214700 $D=9
D49 gnd! OEN dn PJ=0.0002 m=1 $X=31260 $Y=-99700 $D=9
D50 gnd! OEN dn PJ=0.0002 m=1 $X=31260 $Y=110300 $D=9
D51 OEN vdd! dn PJ=0.0002 m=1 $X=33580 $Y=-95300 $D=9
D52 OEN vdd! dn PJ=0.0002 m=1 $X=33580 $Y=114700 $D=9
D53 gnd! OEN dn PJ=0.0002 m=1 $X=35900 $Y=-99700 $D=9
D54 gnd! OEN dn PJ=0.0002 m=1 $X=35900 $Y=110300 $D=9
D55 OEN vdd! dn PJ=0.0002 m=1 $X=38220 $Y=-95300 $D=9
D56 OEN vdd! dn PJ=0.0002 m=1 $X=38220 $Y=114700 $D=9
D57 gnd! OEN dn PJ=0.0001 m=1 $X=40540 $Y=-99700 $D=9
D58 gnd! OEN dn PJ=0.0001 m=1 $X=40540 $Y=110300 $D=9
D59 OEN vdd! dn PJ=0.0001 m=1 $X=43720 $Y=4700 $D=9
D60 OEN vdd! dn PJ=0.0001 m=1 $X=43720 $Y=214700 $D=9
D61 gnd! OEN dn PJ=0.0002 m=1 $X=46040 $Y=-99700 $D=9
D62 gnd! OEN dn PJ=0.0002 m=1 $X=46040 $Y=110300 $D=9
D63 OEN vdd! dn PJ=0.0002 m=1 $X=48360 $Y=-95300 $D=9
D64 OEN vdd! dn PJ=0.0002 m=1 $X=48360 $Y=114700 $D=9
D65 gnd! OEN dn PJ=0.0002 m=1 $X=50680 $Y=-99700 $D=9
D66 gnd! OEN dn PJ=0.0002 m=1 $X=50680 $Y=110300 $D=9
D67 OEN vdd! dn PJ=0.0002 m=1 $X=53000 $Y=-95300 $D=9
D68 OEN vdd! dn PJ=0.0002 m=1 $X=53000 $Y=114700 $D=9
D69 gnd! OEN dn PJ=0.0001 m=1 $X=55320 $Y=-99700 $D=9
D70 gnd! OEN dn PJ=0.0001 m=1 $X=55320 $Y=110300 $D=9
D71 OEN vdd! dn PJ=0.0001 m=1 $X=58500 $Y=4700 $D=9
D72 OEN vdd! dn PJ=0.0001 m=1 $X=58500 $Y=214700 $D=9
D73 gnd! OEN dn PJ=0.0002 m=1 $X=60820 $Y=-99700 $D=9
D74 gnd! OEN dn PJ=0.0002 m=1 $X=60820 $Y=110300 $D=9
D75 OEN vdd! dn PJ=0.0002 m=1 $X=63140 $Y=-95300 $D=9
D76 OEN vdd! dn PJ=0.0002 m=1 $X=63140 $Y=114700 $D=9
D77 gnd! OEN dn PJ=0.0002 m=1 $X=65460 $Y=-99700 $D=9
D78 gnd! OEN dn PJ=0.0002 m=1 $X=65460 $Y=110300 $D=9
D79 OEN vdd! dn PJ=0.0002 m=1 $X=67780 $Y=-95300 $D=9
D80 OEN vdd! dn PJ=0.0002 m=1 $X=67780 $Y=114700 $D=9
D81 gnd! OEN dn PJ=0.0001 m=1 $X=70100 $Y=-99700 $D=9
D82 gnd! OEN dn PJ=0.0001 m=1 $X=70100 $Y=110300 $D=9
D83 OEN vdd! dn PJ=0.0001 m=1 $X=73280 $Y=4700 $D=9
D84 OEN vdd! dn PJ=0.0001 m=1 $X=73280 $Y=214700 $D=9
D85 gnd! OEN dn PJ=0.0002 m=1 $X=75600 $Y=-99700 $D=9
D86 gnd! OEN dn PJ=0.0002 m=1 $X=75600 $Y=110300 $D=9
D87 OEN vdd! dn PJ=0.0002 m=1 $X=77920 $Y=-95300 $D=9
D88 OEN vdd! dn PJ=0.0002 m=1 $X=77920 $Y=114700 $D=9
D89 gnd! OEN dn PJ=0.0002 m=1 $X=80240 $Y=-99700 $D=9
D90 gnd! OEN dn PJ=0.0002 m=1 $X=80240 $Y=110300 $D=9
D91 OEN vdd! dn PJ=0.0002 m=1 $X=82560 $Y=-95300 $D=9
D92 OEN vdd! dn PJ=0.0002 m=1 $X=82560 $Y=114700 $D=9
D93 gnd! OEN dn PJ=0.0001 m=1 $X=84880 $Y=-99700 $D=9
D94 gnd! OEN dn PJ=0.0001 m=1 $X=84880 $Y=110300 $D=9
D95 OEN vdd! dn PJ=0.0001 m=1 $X=88060 $Y=4700 $D=9
D96 OEN vdd! dn PJ=0.0001 m=1 $X=88060 $Y=214700 $D=9
D97 gnd! OEN dn PJ=0.0002 m=1 $X=90380 $Y=-99700 $D=9
D98 gnd! OEN dn PJ=0.0002 m=1 $X=90380 $Y=110300 $D=9
D99 OEN vdd! dn PJ=0.0002 m=1 $X=92700 $Y=-95300 $D=9
D100 OEN vdd! dn PJ=0.0002 m=1 $X=92700 $Y=114700 $D=9
D101 gnd! OEN dn PJ=0.0002 m=1 $X=95020 $Y=-99700 $D=9
D102 gnd! OEN dn PJ=0.0002 m=1 $X=95020 $Y=110300 $D=9
D103 gnd! 17 dn PJ=5e-06 m=1 $X=1560 $Y=328560 $D=10
D104 17 vdd! dn PJ=5e-06 m=1 $X=1560 $Y=334960 $D=10
D105 gnd! 17 dn PJ=5e-06 m=1 $X=1560 $Y=329900 $D=11
D106 17 vdd! dn PJ=5e-06 m=1 $X=1560 $Y=332220 $D=11
X121 gnd! vdd! cpoly_p_CDNS_5887047866511 $T=8060 317780 0 0 $X=8060 $Y=317780
X122 vdd! gnd! cpoly_n_CDNS_5887047866514 $T=540 336500 0 0 $X=540 $Y=336500
X123 OEN 17 PAD $T=0 1440 0 0 $X=-5000 $Y=-235000
X124 vdd! gnd! cpoly_n_CDNS_5887047866566 $T=64300 328000 0 0 $X=64300 $Y=328000
X125 vdd! gnd! cpoly_n_CDNS_5887047866566 $T=73600 328000 0 0 $X=73600 $Y=328000
X126 vdd! gnd! cpoly_n_CDNS_5887047866566 $T=83680 328000 0 0 $X=83680 $Y=328000
X127 gnd! 9 vdd! 8 ICV_87 $T=18620 326300 0 0 $X=18620 $Y=326300
X128 gnd! 9 vdd! 8 ICV_87 $T=23260 326300 0 0 $X=23260 $Y=326300
X129 gnd! nOE_Master vdd! 9 ICV_87 $T=30380 326100 0 0 $X=30380 $Y=326100
X130 gnd! nOE_Master vdd! 9 ICV_87 $T=35020 326100 0 0 $X=35020 $Y=326100
X131 gnd! nOE_Master vdd! 9 ICV_87 $T=39660 326300 0 0 $X=39660 $Y=326300
X132 gnd! nOE_Master vdd! 9 ICV_87 $T=44300 326300 0 0 $X=44300 $Y=326300
X133 gnd! nOE_Master vdd! 9 ICV_87 $T=48940 326300 0 0 $X=48940 $Y=326300
X134 gnd! nOE_Master vdd! 9 ICV_87 $T=53580 326300 0 0 $X=53580 $Y=326300
X135 gnd! nOE_Master vdd! 9 ICV_87 $T=58220 326300 0 0 $X=58220 $Y=326300
X136 gnd! nOE_Master vdd! 9 ICV_87 $T=62860 326300 0 0 $X=62860 $Y=326300
.ENDS
***************************************
.SUBCKT ICV_88 1 2 3 4
** N=4 EP=4 IP=12 FDC=4
M0 2 4 1 1 nmos_a L=2.4e-07 W=2.4e-06 AD=1.4e-12 AS=6.24e-13 PD=3.5e-06 PS=1.75e-06 w_cont=1.1e-06 nfing=1 source_num=2 $X=-140 $Y=200 $D=1
M1 2 4 1 1 nmos_a L=2.4e-07 W=2.4e-06 AD=1.4e-12 AS=6.24e-13 PD=3.5e-06 PS=1.75e-06 w_cont=1.1e-06 nfing=1 source_num=2 $X=620 $Y=200 $D=1
M2 2 4 3 3 pmos_a L=2.4e-07 W=4.5e-06 AD=2.04e-12 AS=1.785e-13 PD=5.1e-06 PS=2.55e-06 w_cont=6e-07 nfing=1 mmm=1 $X=-140 $Y=4600 $D=5
M3 2 4 3 3 pmos_a L=2.4e-07 W=4.5e-06 AD=2.04e-12 AS=1.785e-13 PD=5.1e-06 PS=2.55e-06 w_cont=6e-07 nfing=1 mmm=1 $X=620 $Y=4600 $D=5
.ENDS
***************************************
.SUBCKT PADIN_CE nATD4 nATD3 nATD2 CS nClk gnd! vdd! CEN nATD1 CE
** N=27 EP=10 IP=158 FDC=252
M0 13 11 gnd! gnd! nmos_a L=2.4e-07 W=1.2e-06 AD=7.2e-13 AS=4.8e-13 PD=1.8e-06 PS=9e-07 w_cont=6e-07 nfing=1 source_num=2 $X=19400 $Y=329320 $D=1
M1 13 24 gnd! gnd! nmos_a L=2.4e-07 W=1.2e-06 AD=7.2e-13 AS=4.8e-13 PD=1.8e-06 PS=9e-07 w_cont=6e-07 nfing=1 source_num=2 $X=20840 $Y=329320 $D=1
M2 16 13 gnd! gnd! nmos_a L=2.4e-07 W=2.4e-06 AD=9.1e-13 AS=9.6e-13 PD=1.75e-06 PS=1.75e-06 w_cont=1.1e-06 nfing=1 source_num=2 $X=25540 $Y=326540 $D=1
M3 16 13 gnd! gnd! nmos_a L=2.4e-07 W=2.4e-06 AD=9.1e-13 AS=9.6e-13 PD=1.75e-06 PS=1.75e-06 w_cont=1.1e-06 nfing=1 source_num=2 $X=26300 $Y=326540 $D=1
M4 22 nATD4 19 19 nmos_a L=2.4e-07 W=1.2e-06 AD=7.2e-13 AS=4.8e-13 PD=1.8e-06 PS=9e-07 w_cont=6e-07 nfing=1 source_num=2 $X=12920 $Y=328420 $D=1
M5 19 nATD3 20 20 nmos_a L=2.4e-07 W=1.2e-06 AD=7.2e-13 AS=4.8e-13 PD=1.8e-06 PS=9e-07 w_cont=6e-07 nfing=1 source_num=2 $X=14360 $Y=328420 $D=1
M6 20 nATD2 21 21 nmos_a L=2.4e-07 W=1.2e-06 AD=7.2e-13 AS=4.8e-13 PD=1.8e-06 PS=9e-07 w_cont=6e-07 nfing=1 source_num=2 $X=15800 $Y=328420 $D=1
M7 21 nATD1 gnd! gnd! nmos_a L=2.4e-07 W=1.2e-06 AD=7.2e-13 AS=6.24e-13 PD=1.8e-06 PS=9e-07 w_cont=6e-07 nfing=1 source_num=2 $X=17240 $Y=328740 $D=1
M8 12 22 gnd! gnd! nmos_a L=2.4e-07 W=1.2e-06 AD=7.2e-13 AS=6.24e-13 PD=1.8e-06 PS=9e-07 w_cont=6e-07 nfing=1 source_num=2 $X=18000 $Y=328740 $D=1
M9 17 27 gnd! gnd! nmos_a L=2.4e-07 W=4.8e-07 AD=4.32e-13 AS=1.92e-13 PD=1.08e-06 PS=5.4e-07 w_cont=6e-07 nfing=1 source_num=2 $X=8820 $Y=327700 $D=1
M10 11 17 gnd! gnd! nmos_a L=2.4e-07 W=4.8e-07 AD=4.32e-13 AS=1.92e-13 PD=1.08e-06 PS=5.4e-07 w_cont=6e-07 nfing=1 source_num=2 $X=10260 $Y=327700 $D=1
M11 24 CS gnd! gnd! nmos_a L=2.4e-07 W=4.8e-07 AD=4.32e-13 AS=1.92e-13 PD=1.08e-06 PS=5.4e-07 w_cont=6e-07 nfing=1 source_num=2 $X=22280 $Y=330040 $D=1
M12 25 12 gnd! gnd! nmos_a L=2.4e-07 W=3.6e-06 AD=1.664e-12 AS=1.44e-12 PD=4.16e-06 PS=2.08e-06 w_cont=1.6e-06 nfing=1 source_num=2 $X=27780 $Y=326540 $D=1
M13 26 CE 25 25 nmos_a L=2.4e-07 W=3.6e-06 AD=1.664e-12 AS=1.44e-12 PD=4.16e-06 PS=2.08e-06 w_cont=1.6e-06 nfing=1 source_num=2 $X=29220 $Y=326540 $D=1
M14 14 13 26 26 nmos_a L=2.4e-07 W=3.6e-06 AD=1.664e-12 AS=1.44e-12 PD=4.16e-06 PS=2.08e-06 w_cont=1.6e-06 nfing=1 source_num=2 $X=30660 $Y=326540 $D=1
M15 18 11 vdd! vdd! pmos_a L=4e-07 W=4.8e-07 AD=4.32e-13 AS=1.224e-13 PD=1.08e-06 PS=5.4e-07 w_cont=6e-07 nfing=1 mmm=1 $X=10220 $Y=332940 $D=5
M16 13 11 23 23 pmos_a L=2.4e-07 W=2.88e-06 AD=1.392e-12 AS=1.344e-13 PD=3.48e-06 PS=1.74e-06 w_cont=6e-07 nfing=1 mmm=1 $X=19400 $Y=332000 $D=5
M17 23 24 vdd! vdd! pmos_a L=2.4e-07 W=2.88e-06 AD=1.392e-12 AS=1.344e-13 PD=3.48e-06 PS=1.74e-06 w_cont=6e-07 nfing=1 mmm=1 $X=20840 $Y=332000 $D=5
M18 14 12 vdd! vdd! pmos_a L=2.4e-07 W=2.22e-06 AD=1.128e-12 AS=1.311e-13 PD=2.82e-06 PS=1.41e-06 w_cont=6e-07 nfing=1 mmm=1 $X=27780 $Y=332660 $D=5
M19 14 CE vdd! vdd! pmos_a L=2.4e-07 W=2.22e-06 AD=1.128e-12 AS=1.311e-13 PD=2.82e-06 PS=1.41e-06 w_cont=6e-07 nfing=1 mmm=1 $X=29220 $Y=332660 $D=5
M20 14 13 vdd! vdd! pmos_a L=2.4e-07 W=2.22e-06 AD=1.128e-12 AS=1.311e-13 PD=2.82e-06 PS=1.41e-06 w_cont=6e-07 nfing=1 mmm=1 $X=30660 $Y=332660 $D=5
M21 12 22 vdd! vdd! pmos_a L=2.4e-07 W=2e-06 AD=1.04e-12 AS=1.3e-13 PD=2.6e-06 PS=1.3e-06 w_cont=6e-07 nfing=1 mmm=1 $X=18000 $Y=331860 $D=5
M22 18 27 vdd! vdd! pmos_a L=2.4e-07 W=1e-06 AD=6.4e-13 AS=1.25e-13 PD=1.6e-06 PS=8e-07 w_cont=6e-07 nfing=1 mmm=1 $X=8820 $Y=332940 $D=5
M23 17 27 18 18 pmos_a L=2.4e-07 W=1e-06 AD=6.4e-13 AS=1.25e-13 PD=1.6e-06 PS=8e-07 w_cont=6e-07 nfing=1 mmm=1 $X=8820 $Y=330300 $D=5
M24 11 17 vdd! vdd! pmos_a L=2.4e-07 W=1e-06 AD=6.4e-13 AS=1.25e-13 PD=1.6e-06 PS=8e-07 w_cont=6e-07 nfing=1 mmm=1 $X=10260 $Y=330140 $D=5
M25 22 nATD4 vdd! vdd! pmos_a L=2.4e-07 W=1e-06 AD=6.4e-13 AS=1.25e-13 PD=1.6e-06 PS=8e-07 w_cont=6e-07 nfing=1 mmm=1 $X=12920 $Y=332860 $D=5
M26 22 nATD3 vdd! vdd! pmos_a L=2.4e-07 W=1e-06 AD=6.4e-13 AS=1.61e-13 PD=1.6e-06 PS=8e-07 w_cont=6e-07 nfing=1 mmm=1 $X=14360 $Y=332860 $D=5
M27 22 nATD2 vdd! vdd! pmos_a L=2.4e-07 W=1e-06 AD=6.4e-13 AS=1.61e-13 PD=1.6e-06 PS=8e-07 w_cont=6e-07 nfing=1 mmm=1 $X=15120 $Y=332860 $D=5
M28 22 nATD1 vdd! vdd! pmos_a L=2.4e-07 W=1e-06 AD=6.4e-13 AS=1.25e-13 PD=1.6e-06 PS=8e-07 w_cont=6e-07 nfing=1 mmm=1 $X=16560 $Y=332860 $D=5
M29 24 CS vdd! vdd! pmos_a L=2.4e-07 W=1e-06 AD=6.4e-13 AS=1.25e-13 PD=1.6e-06 PS=8e-07 w_cont=6e-07 nfing=1 mmm=1 $X=22280 $Y=332500 $D=5
M30 16 13 vdd! vdd! pmos_a L=2.4e-07 W=4e-06 AD=1.84e-12 AS=1.76e-13 PD=4.6e-06 PS=2.3e-06 w_cont=6e-07 nfing=1 mmm=1 $X=25540 $Y=330880 $D=5
M31 16 13 vdd! vdd! pmos_a L=2.4e-07 W=4e-06 AD=1.84e-12 AS=1.76e-13 PD=4.6e-06 PS=2.3e-06 w_cont=6e-07 nfing=1 mmm=1 $X=26300 $Y=330880 $D=5
M32 vdd! gnd! vdd! cpoly_n w=6e-06 l=2e-06 c=7.5402e-14 as=2.4e-13 ad=2.304e-12 ps=2.88e-06 pd=4.86761e-06 sim_w=5.76e-06 m_per_maxw=1.04167 numb_sub_cont=3 nfing=1 $X=34260 $Y=328200 $D=22
M33 vdd! gnd! vdd! cpoly_n w=6e-06 l=2e-06 c=7.5402e-14 as=2.4e-13 ad=2.304e-12 ps=2.88e-06 pd=4.86761e-06 sim_w=5.76e-06 m_per_maxw=1.04167 numb_sub_cont=3 nfing=1 $X=39620 $Y=328200 $D=22
M34 vdd! gnd! vdd! cpoly_n w=6e-06 l=2e-06 c=7.5402e-14 as=2.4e-13 ad=2.304e-12 ps=2.88e-06 pd=4.86761e-06 sim_w=5.76e-06 m_per_maxw=1.04167 numb_sub_cont=3 nfing=1 $X=45020 $Y=328200 $D=22
M35 vdd! gnd! vdd! cpoly_n w=6e-06 l=2e-06 c=7.5402e-14 as=2.4e-13 ad=2.304e-12 ps=2.88e-06 pd=4.86761e-06 sim_w=5.76e-06 m_per_maxw=1.04167 numb_sub_cont=3 nfing=1 $X=50420 $Y=328200 $D=22
M36 vdd! gnd! vdd! cpoly_n w=6e-06 l=2e-06 c=7.5402e-14 as=2.4e-13 ad=2.304e-12 ps=2.88e-06 pd=4.86761e-06 sim_w=5.76e-06 m_per_maxw=1.04167 numb_sub_cont=3 nfing=1 $X=55820 $Y=328200 $D=22
M37 vdd! gnd! vdd! cpoly_n w=6e-06 l=2e-06 c=7.5402e-14 as=2.4e-13 ad=2.304e-12 ps=2.88e-06 pd=4.86761e-06 sim_w=5.76e-06 m_per_maxw=1.04167 numb_sub_cont=3 nfing=1 $X=61220 $Y=328200 $D=22
M38 vdd! gnd! vdd! cpoly_n w=6e-06 l=2e-06 c=7.5402e-14 as=2.4e-13 ad=2.304e-12 ps=2.88e-06 pd=4.86761e-06 sim_w=5.76e-06 m_per_maxw=1.04167 numb_sub_cont=3 nfing=1 $X=66600 $Y=328200 $D=22
M39 vdd! gnd! vdd! cpoly_n w=6e-06 l=2e-06 c=7.5402e-14 as=2.4e-13 ad=2.304e-12 ps=2.88e-06 pd=4.86761e-06 sim_w=5.76e-06 m_per_maxw=1.04167 numb_sub_cont=3 nfing=1 $X=71960 $Y=328200 $D=22
M40 vdd! gnd! vdd! cpoly_n w=6e-06 l=2e-06 c=7.5402e-14 as=2.4e-13 ad=2.304e-12 ps=2.88e-06 pd=4.86761e-06 sim_w=5.76e-06 m_per_maxw=1.04167 numb_sub_cont=3 nfing=1 $X=77320 $Y=328200 $D=22
M41 vdd! gnd! vdd! cpoly_n w=6e-06 l=2e-06 c=7.5402e-14 as=2.4e-13 ad=2.304e-12 ps=2.88e-06 pd=4.86761e-06 sim_w=5.76e-06 m_per_maxw=1.04167 numb_sub_cont=3 nfing=1 $X=82720 $Y=328200 $D=22
M42 vdd! gnd! vdd! cpoly_n w=6e-06 l=2e-06 c=7.5402e-14 as=2.4e-13 ad=2.304e-12 ps=2.88e-06 pd=4.86761e-06 sim_w=5.76e-06 m_per_maxw=1.04167 numb_sub_cont=3 nfing=1 $X=88120 $Y=328200 $D=22
M43 vdd! gnd! vdd! cpoly_n w=6e-06 l=2e-06 c=7.5402e-14 as=2.4e-13 ad=2.304e-12 ps=2.88e-06 pd=4.86761e-06 sim_w=5.76e-06 m_per_maxw=1.04167 numb_sub_cont=3 nfing=1 $X=93520 $Y=328200 $D=22
D44 CEN vdd! dn PJ=0.0002 m=1 $X=4020 $Y=-95300 $D=9
D45 CEN vdd! dn PJ=0.0002 m=1 $X=4020 $Y=114700 $D=9
D46 gnd! CEN dn PJ=0.0002 m=1 $X=6340 $Y=-99700 $D=9
D47 gnd! CEN dn PJ=0.0002 m=1 $X=6340 $Y=110300 $D=9
D48 CEN vdd! dn PJ=0.0002 m=1 $X=8660 $Y=-95300 $D=9
D49 CEN vdd! dn PJ=0.0002 m=1 $X=8660 $Y=114700 $D=9
D50 gnd! CEN dn PJ=0.0001 m=1 $X=10980 $Y=-99700 $D=9
D51 gnd! CEN dn PJ=0.0001 m=1 $X=10980 $Y=110300 $D=9
D52 CEN vdd! dn PJ=0.0001 m=1 $X=14160 $Y=4700 $D=9
D53 CEN vdd! dn PJ=0.0001 m=1 $X=14160 $Y=214700 $D=9
D54 gnd! CEN dn PJ=0.0002 m=1 $X=16480 $Y=-99700 $D=9
D55 gnd! CEN dn PJ=0.0002 m=1 $X=16480 $Y=110300 $D=9
D56 CEN vdd! dn PJ=0.0002 m=1 $X=18800 $Y=-95300 $D=9
D57 CEN vdd! dn PJ=0.0002 m=1 $X=18800 $Y=114700 $D=9
D58 gnd! CEN dn PJ=0.0002 m=1 $X=21120 $Y=-99700 $D=9
D59 gnd! CEN dn PJ=0.0002 m=1 $X=21120 $Y=110300 $D=9
D60 CEN vdd! dn PJ=0.0002 m=1 $X=23440 $Y=-95300 $D=9
D61 CEN vdd! dn PJ=0.0002 m=1 $X=23440 $Y=114700 $D=9
D62 gnd! CEN dn PJ=0.0001 m=1 $X=25760 $Y=-99700 $D=9
D63 gnd! CEN dn PJ=0.0001 m=1 $X=25760 $Y=110300 $D=9
D64 CEN vdd! dn PJ=0.0001 m=1 $X=28940 $Y=4700 $D=9
D65 CEN vdd! dn PJ=0.0001 m=1 $X=28940 $Y=214700 $D=9
D66 gnd! CEN dn PJ=0.0002 m=1 $X=31260 $Y=-99700 $D=9
D67 gnd! CEN dn PJ=0.0002 m=1 $X=31260 $Y=110300 $D=9
D68 CEN vdd! dn PJ=0.0002 m=1 $X=33580 $Y=-95300 $D=9
D69 CEN vdd! dn PJ=0.0002 m=1 $X=33580 $Y=114700 $D=9
D70 gnd! CEN dn PJ=0.0002 m=1 $X=35900 $Y=-99700 $D=9
D71 gnd! CEN dn PJ=0.0002 m=1 $X=35900 $Y=110300 $D=9
D72 CEN vdd! dn PJ=0.0002 m=1 $X=38220 $Y=-95300 $D=9
D73 CEN vdd! dn PJ=0.0002 m=1 $X=38220 $Y=114700 $D=9
D74 gnd! CEN dn PJ=0.0001 m=1 $X=40540 $Y=-99700 $D=9
D75 gnd! CEN dn PJ=0.0001 m=1 $X=40540 $Y=110300 $D=9
D76 CEN vdd! dn PJ=0.0001 m=1 $X=43720 $Y=4700 $D=9
D77 CEN vdd! dn PJ=0.0001 m=1 $X=43720 $Y=214700 $D=9
D78 gnd! CEN dn PJ=0.0002 m=1 $X=46040 $Y=-99700 $D=9
D79 gnd! CEN dn PJ=0.0002 m=1 $X=46040 $Y=110300 $D=9
D80 CEN vdd! dn PJ=0.0002 m=1 $X=48360 $Y=-95300 $D=9
D81 CEN vdd! dn PJ=0.0002 m=1 $X=48360 $Y=114700 $D=9
D82 gnd! CEN dn PJ=0.0002 m=1 $X=50680 $Y=-99700 $D=9
D83 gnd! CEN dn PJ=0.0002 m=1 $X=50680 $Y=110300 $D=9
D84 CEN vdd! dn PJ=0.0002 m=1 $X=53000 $Y=-95300 $D=9
D85 CEN vdd! dn PJ=0.0002 m=1 $X=53000 $Y=114700 $D=9
D86 gnd! CEN dn PJ=0.0001 m=1 $X=55320 $Y=-99700 $D=9
D87 gnd! CEN dn PJ=0.0001 m=1 $X=55320 $Y=110300 $D=9
D88 CEN vdd! dn PJ=0.0001 m=1 $X=58500 $Y=4700 $D=9
D89 CEN vdd! dn PJ=0.0001 m=1 $X=58500 $Y=214700 $D=9
D90 gnd! CEN dn PJ=0.0002 m=1 $X=60820 $Y=-99700 $D=9
D91 gnd! CEN dn PJ=0.0002 m=1 $X=60820 $Y=110300 $D=9
D92 CEN vdd! dn PJ=0.0002 m=1 $X=63140 $Y=-95300 $D=9
D93 CEN vdd! dn PJ=0.0002 m=1 $X=63140 $Y=114700 $D=9
D94 gnd! CEN dn PJ=0.0002 m=1 $X=65460 $Y=-99700 $D=9
D95 gnd! CEN dn PJ=0.0002 m=1 $X=65460 $Y=110300 $D=9
D96 CEN vdd! dn PJ=0.0002 m=1 $X=67780 $Y=-95300 $D=9
D97 CEN vdd! dn PJ=0.0002 m=1 $X=67780 $Y=114700 $D=9
D98 gnd! CEN dn PJ=0.0001 m=1 $X=70100 $Y=-99700 $D=9
D99 gnd! CEN dn PJ=0.0001 m=1 $X=70100 $Y=110300 $D=9
D100 CEN vdd! dn PJ=0.0001 m=1 $X=73280 $Y=4700 $D=9
D101 CEN vdd! dn PJ=0.0001 m=1 $X=73280 $Y=214700 $D=9
D102 gnd! CEN dn PJ=0.0002 m=1 $X=75600 $Y=-99700 $D=9
D103 gnd! CEN dn PJ=0.0002 m=1 $X=75600 $Y=110300 $D=9
D104 CEN vdd! dn PJ=0.0002 m=1 $X=77920 $Y=-95300 $D=9
D105 CEN vdd! dn PJ=0.0002 m=1 $X=77920 $Y=114700 $D=9
D106 gnd! CEN dn PJ=0.0002 m=1 $X=80240 $Y=-99700 $D=9
D107 gnd! CEN dn PJ=0.0002 m=1 $X=80240 $Y=110300 $D=9
D108 CEN vdd! dn PJ=0.0002 m=1 $X=82560 $Y=-95300 $D=9
D109 CEN vdd! dn PJ=0.0002 m=1 $X=82560 $Y=114700 $D=9
D110 gnd! CEN dn PJ=0.0001 m=1 $X=84880 $Y=-99700 $D=9
D111 gnd! CEN dn PJ=0.0001 m=1 $X=84880 $Y=110300 $D=9
D112 CEN vdd! dn PJ=0.0001 m=1 $X=88060 $Y=4700 $D=9
D113 CEN vdd! dn PJ=0.0001 m=1 $X=88060 $Y=214700 $D=9
D114 gnd! CEN dn PJ=0.0002 m=1 $X=90380 $Y=-99700 $D=9
D115 gnd! CEN dn PJ=0.0002 m=1 $X=90380 $Y=110300 $D=9
D116 CEN vdd! dn PJ=0.0002 m=1 $X=92700 $Y=-95300 $D=9
D117 CEN vdd! dn PJ=0.0002 m=1 $X=92700 $Y=114700 $D=9
D118 gnd! CEN dn PJ=0.0002 m=1 $X=95020 $Y=-99700 $D=9
D119 gnd! CEN dn PJ=0.0002 m=1 $X=95020 $Y=110300 $D=9
D120 gnd! 27 dn PJ=5e-06 m=1 $X=1560 $Y=328560 $D=10
D121 27 vdd! dn PJ=5e-06 m=1 $X=1560 $Y=334960 $D=10
D122 gnd! 27 dn PJ=5e-06 m=1 $X=1560 $Y=329900 $D=11
D123 27 vdd! dn PJ=5e-06 m=1 $X=1560 $Y=332220 $D=11
X158 gnd! vdd! cpoly_p_CDNS_5887047866511 $T=7840 317780 0 0 $X=7840 $Y=317780
X159 vdd! gnd! cpoly_n_CDNS_5887047866514 $T=520 336500 0 0 $X=520 $Y=336500
X160 CEN 27 PAD $T=0 1440 0 0 $X=-5000 $Y=-235000
X163 gnd! 15 vdd! 14 ICV_88 $T=32920 326300 1 180 $X=31480 $Y=326300
X164 gnd! 15 vdd! 14 ICV_88 $T=38280 326300 1 180 $X=36840 $Y=326300
X165 gnd! nClk vdd! 15 ICV_88 $T=43680 326300 1 180 $X=42240 $Y=326300
X166 gnd! nClk vdd! 15 ICV_88 $T=49080 326300 1 180 $X=47640 $Y=326300
X167 gnd! nClk vdd! 15 ICV_88 $T=54480 326300 1 180 $X=53040 $Y=326300
X168 gnd! nClk vdd! 15 ICV_88 $T=59880 326300 1 180 $X=58440 $Y=326300
X169 gnd! nClk vdd! 15 ICV_88 $T=65260 326300 1 180 $X=63820 $Y=326300
X170 gnd! nClk vdd! 15 ICV_88 $T=70620 326300 1 180 $X=69180 $Y=326300
X171 gnd! nClk vdd! 15 ICV_88 $T=75980 326100 1 180 $X=74540 $Y=326100
X172 gnd! CE vdd! 16 ICV_88 $T=81380 326080 1 180 $X=79940 $Y=326080
X173 gnd! CE vdd! 16 ICV_88 $T=86780 326080 1 180 $X=85340 $Y=326080
X174 gnd! CE vdd! 16 ICV_88 $T=92180 326080 1 180 $X=90740 $Y=326080
X175 gnd! CE vdd! 16 ICV_88 $T=97580 326080 1 180 $X=96140 $Y=326080
.ENDS
***************************************
.SUBCKT nmos_a_CDNS_5887047866520 1 2 3
** N=3 EP=3 IP=0 FDC=1
M0 2 3 1 1 nmos_a L=2.4e-07 W=1e-06 AD=6.4e-13 AS=4e-13 PD=1.6e-06 PS=8e-07 w_cont=6e-07 nfing=1 source_num=2 $X=620 $Y=200 $D=1
.ENDS
***************************************
.SUBCKT PADIN_CS gnd! vdd! CS nE nCS
** N=13 EP=5 IP=104 FDC=129
M0 8 11 vdd! vdd! pmos_a L=4e-07 W=4.8e-07 AD=5.71272e-13 AS=1.224e-13 PD=4.35224e-07 PS=5.4e-07 w_cont=6e-07 nfing=1 mmm=1 $X=10520 $Y=333300 $D=5
M1 11 10 vdd! vdd! pmos_a L=2.4e-07 W=1e-06 AD=6.4e-13 AS=1.25e-13 PD=1.6e-06 PS=8e-07 w_cont=6e-07 nfing=1 mmm=1 $X=12160 $Y=332780 $D=5
M2 6 11 vdd! vdd! pmos_a L=2.4e-07 W=2e-06 AD=1.04e-12 AS=1.3e-13 PD=2.6e-06 PS=1.3e-06 w_cont=6e-07 nfing=1 mmm=1 $X=13600 $Y=331520 $D=5
M3 8 8 vdd! vdd! pmos_a L=2.4e-07 W=1e-06 AD=8.46328e-13 AS=1.25e-13 PD=9.55224e-07 PS=8e-07 w_cont=6e-07 nfing=1 mmm=1 $X=9160 $Y=332980 $D=5
M4 10 13 8 8 pmos_a L=2.4e-07 W=1e-06 AD=6.4e-13 AS=1.25e-13 PD=1.6e-06 PS=8e-07 w_cont=6e-07 nfing=1 mmm=1 $X=9240 $Y=330180 $D=5
M5 12 nE vdd! vdd! pmos_a L=2.4e-07 W=1e-06 AD=6.4e-13 AS=1.25e-13 PD=1.6e-06 PS=8e-07 w_cont=6e-07 nfing=1 mmm=1 $X=15000 $Y=331520 $D=5
M6 10 12 vdd! vdd! pmos_a L=2.4e-07 W=4.8e-07 AD=4.32e-13 AS=1.224e-13 PD=1.08e-06 PS=5.4e-07 w_cont=6e-07 nfing=1 mmm=1 $X=10680 $Y=330180 $D=5
M7 vdd! gnd! vdd! cpoly_n w=6e-06 l=2e-06 c=7.5402e-14 as=2.4e-13 ad=2.304e-12 ps=2.88e-06 pd=4.86761e-06 sim_w=5.76e-06 m_per_maxw=1.04167 numb_sub_cont=3 nfing=1 $X=20680 $Y=328200 $D=22
M8 vdd! gnd! vdd! cpoly_n w=6e-06 l=2e-06 c=7.5402e-14 as=3.0336e-13 ad=2.304e-12 ps=2.88e-06 pd=4.86761e-06 sim_w=5.76e-06 m_per_maxw=1.04167 numb_sub_cont=3 nfing=1 $X=25280 $Y=328200 $D=22
M9 vdd! gnd! vdd! cpoly_n w=6e-06 l=2e-06 c=7.5402e-14 as=3.0336e-13 ad=2.304e-12 ps=2.88e-06 pd=4.86761e-06 sim_w=5.76e-06 m_per_maxw=1.04167 numb_sub_cont=3 nfing=1 $X=27800 $Y=328200 $D=22
M10 vdd! gnd! vdd! cpoly_n w=6e-06 l=2e-06 c=7.5402e-14 as=2.4e-13 ad=2.304e-12 ps=2.88e-06 pd=4.86761e-06 sim_w=5.76e-06 m_per_maxw=1.04167 numb_sub_cont=3 nfing=1 $X=32440 $Y=328200 $D=22
M11 vdd! gnd! vdd! cpoly_n w=6e-06 l=2e-06 c=7.5402e-14 as=2.4e-13 ad=2.304e-12 ps=2.88e-06 pd=4.86761e-06 sim_w=5.76e-06 m_per_maxw=1.04167 numb_sub_cont=3 nfing=1 $X=37080 $Y=328200 $D=22
M12 vdd! gnd! vdd! cpoly_n w=6e-06 l=2e-06 c=7.5402e-14 as=2.4e-13 ad=2.304e-12 ps=2.88e-06 pd=4.86761e-06 sim_w=5.76e-06 m_per_maxw=1.04167 numb_sub_cont=3 nfing=1 $X=41720 $Y=328200 $D=22
M13 vdd! gnd! vdd! cpoly_n w=6e-06 l=2e-06 c=7.5402e-14 as=2.4e-13 ad=2.304e-12 ps=2.88e-06 pd=4.86761e-06 sim_w=5.76e-06 m_per_maxw=1.04167 numb_sub_cont=3 nfing=1 $X=46360 $Y=328200 $D=22
M14 vdd! gnd! vdd! cpoly_n w=6e-06 l=2e-06 c=7.5402e-14 as=2.4e-13 ad=2.304e-12 ps=2.88e-06 pd=4.86761e-06 sim_w=5.76e-06 m_per_maxw=1.04167 numb_sub_cont=3 nfing=1 $X=51000 $Y=328200 $D=22
M15 vdd! gnd! vdd! cpoly_n w=6e-06 l=2e-06 c=7.5402e-14 as=2.4e-13 ad=2.304e-12 ps=2.88e-06 pd=4.86761e-06 sim_w=5.76e-06 m_per_maxw=1.04167 numb_sub_cont=3 nfing=1 $X=55640 $Y=328200 $D=22
M16 vdd! gnd! vdd! cpoly_n w=6e-06 l=2e-06 c=7.5402e-14 as=2.4e-13 ad=2.304e-12 ps=2.88e-06 pd=4.86761e-06 sim_w=5.76e-06 m_per_maxw=1.04167 numb_sub_cont=3 nfing=1 $X=60280 $Y=328200 $D=22
M17 vdd! gnd! vdd! cpoly_n w=6e-06 l=2e-06 c=7.5402e-14 as=2.4e-13 ad=2.304e-12 ps=2.88e-06 pd=4.86761e-06 sim_w=5.76e-06 m_per_maxw=1.04167 numb_sub_cont=3 nfing=1 $X=64920 $Y=328200 $D=22
D18 gnd! 13 dn PJ=5e-06 m=1 $X=1560 $Y=328560 $D=10
D19 13 vdd! dn PJ=5e-06 m=1 $X=1560 $Y=334960 $D=10
D20 gnd! 13 dn PJ=5e-06 m=1 $X=1560 $Y=329900 $D=11
D21 13 vdd! dn PJ=5e-06 m=1 $X=1560 $Y=332220 $D=11
X38 gnd! vdd! cpoly_p_CDNS_5887047866511 $T=8060 317780 0 0 $X=8060 $Y=317780
X39 vdd! gnd! cpoly_n_CDNS_5887047866514 $T=540 336500 0 0 $X=540 $Y=336500
X40 CS 13 PAD $T=0 1440 0 0 $X=-5000 $Y=-235000
X41 vdd! gnd! cpoly_n_CDNS_5887047866515 $T=97780 328000 1 180 $X=81940 $Y=328000
X42 gnd! 11 10 nmos_a_CDNS_5887047866521 $T=11540 327980 0 0 $X=11540 $Y=327980
X43 gnd! 12 nE nmos_a_CDNS_5887047866521 $T=15860 329980 0 180 $X=14420 $Y=328480
X44 gnd! 7 vdd! 6 ICV_87 $T=18620 326300 0 0 $X=18620 $Y=326300
X45 gnd! 7 vdd! 6 ICV_87 $T=23260 326300 0 0 $X=23260 $Y=326300
X46 gnd! nCS vdd! 7 ICV_87 $T=30380 326100 0 0 $X=30380 $Y=326100
X47 gnd! nCS vdd! 7 ICV_87 $T=35020 326100 0 0 $X=35020 $Y=326100
X48 gnd! nCS vdd! 7 ICV_87 $T=39660 326300 0 0 $X=39660 $Y=326300
X49 gnd! nCS vdd! 7 ICV_87 $T=44300 326300 0 0 $X=44300 $Y=326300
X50 gnd! nCS vdd! 7 ICV_87 $T=48940 326300 0 0 $X=48940 $Y=326300
X51 gnd! nCS vdd! 7 ICV_87 $T=53580 326300 0 0 $X=53580 $Y=326300
X52 gnd! nCS vdd! 7 ICV_87 $T=58220 326300 0 0 $X=58220 $Y=326300
X53 gnd! nCS vdd! 7 ICV_87 $T=62860 326300 0 0 $X=62860 $Y=326300
X54 9 10 13 nmos_a_CDNS_5887047866520 $T=10100 327480 1 180 $X=8660 $Y=327480
X55 gnd! 9 12 nmos_a_CDNS_5887047866520 $T=11540 327480 1 180 $X=10100 $Y=327480
X56 gnd! 6 11 nmos_a_CDNS_5887047866520 $T=12980 327980 0 0 $X=12980 $Y=327980
.ENDS
***************************************
.SUBCKT nmos_a_CDNS_5887047866581
** N=3 EP=0 IP=0 FDC=0
*.SEEDPROM
.ENDS
***************************************
.SUBCKT pmos_a_CDNS_5887047866583
** N=3 EP=0 IP=0 FDC=0
*.SEEDPROM
.ENDS
***************************************
.SUBCKT pmos_a_CDNS_5887047866580 1 2 3
** N=3 EP=3 IP=0 FDC=1
*.SEEDPROM
M0 2 3 1 1 pmos_a L=2.4e-07 W=2.4e-06 AD=7.8e-13 AS=1.32e-13 PD=1.5e-06 PS=1.5e-06 w_cont=6e-07 nfing=1 mmm=1 $X=620 $Y=200 $D=5
.ENDS
***************************************
.SUBCKT RingPad_EOR In2 In1 Out gnd! vdd! 10
** N=10 EP=6 IP=33 FDC=20
*.SEEDPROM
M0 6 In2 gnd! gnd! nmos_a L=2.4e-07 W=1.2e-06 AD=7.2e-13 AS=4.8e-13 PD=1.8e-06 PS=9e-07 w_cont=6e-07 nfing=1 source_num=2 $X=-2100 $Y=-3020 $D=1
M1 7 In1 6 6 nmos_a L=2.4e-07 W=1.2e-06 AD=7.2e-13 AS=4.8e-13 PD=1.8e-06 PS=9e-07 w_cont=6e-07 nfing=1 source_num=2 $X=-660 $Y=-3020 $D=1
M2 10 7 8 8 nmos_a L=2.4e-07 W=1.2e-06 AD=4.68e-13 AS=4.8e-13 PD=9e-07 PS=9e-07 w_cont=6e-07 nfing=1 source_num=2 $X=780 $Y=-3020 $D=1
M3 10 7 8 8 nmos_a L=2.4e-07 W=1.2e-06 AD=4.68e-13 AS=4.8e-13 PD=9e-07 PS=9e-07 w_cont=6e-07 nfing=1 source_num=2 $X=1540 $Y=-3020 $D=1
M4 8 In2 gnd! gnd! nmos_a L=2.4e-07 W=1.2e-06 AD=4.68e-13 AS=4.8e-13 PD=9e-07 PS=9e-07 w_cont=6e-07 nfing=1 source_num=2 $X=3020 $Y=-3540 $D=1
M5 8 In2 gnd! gnd! nmos_a L=2.4e-07 W=1.2e-06 AD=4.68e-13 AS=6.24e-13 PD=9e-07 PS=9e-07 w_cont=6e-07 nfing=1 source_num=2 $X=3780 $Y=-3540 $D=1
M6 8 In1 gnd! gnd! nmos_a L=2.4e-07 W=1.2e-06 AD=4.68e-13 AS=6.24e-13 PD=9e-07 PS=9e-07 w_cont=6e-07 nfing=1 source_num=2 $X=4540 $Y=-3540 $D=1
M7 8 In1 gnd! gnd! nmos_a L=2.4e-07 W=1.2e-06 AD=4.68e-13 AS=4.8e-13 PD=9e-07 PS=9e-07 w_cont=6e-07 nfing=1 source_num=2 $X=5300 $Y=-3540 $D=1
M8 Out 10 vdd! vdd! pmos_a L=2.4e-07 W=2.4e-06 AD=7.8e-13 AS=1.68e-13 PD=1.5e-06 PS=1.5e-06 w_cont=6e-07 nfing=1 mmm=1 $X=5980 $Y=220 $D=5
M9 Out 10 vdd! vdd! pmos_a L=2.4e-07 W=2.4e-06 AD=7.8e-13 AS=1.68e-13 PD=1.5e-06 PS=1.5e-06 w_cont=6e-07 nfing=1 mmm=1 $X=6740 $Y=220 $D=5
M10 Out 10 vdd! vdd! pmos_a L=2.4e-07 W=2.4e-06 AD=7.8e-13 AS=1.68e-13 PD=1.5e-06 PS=1.5e-06 w_cont=6e-07 nfing=1 mmm=1 $X=7500 $Y=220 $D=5
M11 10 7 vdd! vdd! pmos_a L=2.4e-07 W=2.4e-06 AD=1.2e-12 AS=1.32e-13 PD=3e-06 PS=1.5e-06 w_cont=6e-07 nfing=1 mmm=1 $X=780 $Y=-280 $D=5
M12 10 In2 9 9 pmos_a L=2.4e-07 W=2.4e-06 AD=7.8e-13 AS=1.32e-13 PD=1.5e-06 PS=1.5e-06 w_cont=6e-07 nfing=1 mmm=1 $X=2980 $Y=-280 $D=5
M13 9 In1 vdd! vdd! pmos_a L=2.4e-07 W=2.4e-06 AD=7.8e-13 AS=1.68e-13 PD=1.5e-06 PS=1.5e-06 w_cont=6e-07 nfing=1 mmm=1 $X=5220 $Y=220 $D=5
X14 vdd! 7 In2 pmos_a_CDNS_5887047866540 $T=-2720 720 0 0 $X=-2720 $Y=720
X15 vdd! 7 In1 pmos_a_CDNS_5887047866540 $T=-1280 720 0 0 $X=-1280 $Y=720
X18 gnd! Out 10 nmos_a_CDNS_5887047866573 $T=6880 -4380 0 0 $X=6880 $Y=-4380
X23 9 10 In2 pmos_a_CDNS_5887047866580 $T=1600 -480 0 0 $X=1600 $Y=-480
X24 vdd! 9 In1 pmos_a_CDNS_5887047866580 $T=3840 20 0 0 $X=3840 $Y=20
.ENDS
***************************************
.SUBCKT ICV_89
** N=3 EP=0 IP=6 FDC=0
.ENDS
***************************************
.SUBCKT ICV_90
** N=3 EP=0 IP=6 FDC=0
.ENDS
***************************************
.SUBCKT VDD_Core_PAD vdd! gnd!
** N=8 EP=2 IP=21 FDC=78
*.CALIBRE ISOLATED NETS: VDD_PAD!
X0 vdd! gnd! cpoly_n_CDNS_588704786651 $T=520 333340 0 0 $X=520 $Y=333340
X1 gnd! vdd! cpoly_p_CDNS_588704786650 $T=520 320500 0 0 $X=520 $Y=320500
.ENDS
***************************************
.SUBCKT RingPad_Buffer In Out vdd! gnd!
** N=5 EP=4 IP=30 FDC=20
X0 vdd! 5 In pmos_a_CDNS_5887047866574 $T=600 -520 1 90 $X=600 $Y=-520
X1 vdd! Out 5 pmos_a_CDNS_5887047866574 $T=11340 -520 0 90 $X=6340 $Y=-520
X2 vdd! Out 5 pmos_a_CDNS_5887047866574 $T=17480 -520 0 90 $X=12480 $Y=-520
X3 vdd! Out 5 pmos_a_CDNS_5887047866574 $T=23620 -520 0 90 $X=18620 $Y=-520
X4 vdd! Out 5 pmos_a_CDNS_5887047866574 $T=29760 -520 0 90 $X=24760 $Y=-520
X5 gnd! 5 In nmos_a_CDNS_5887047866573 $T=1200 1720 1 90 $X=1200 $Y=1720
X6 gnd! Out 5 nmos_a_CDNS_5887047866573 $T=10740 1720 0 90 $X=6840 $Y=1720
X7 gnd! Out 5 nmos_a_CDNS_5887047866573 $T=16880 1720 0 90 $X=12980 $Y=1720
X8 gnd! Out 5 nmos_a_CDNS_5887047866573 $T=23020 1720 0 90 $X=19120 $Y=1720
X9 gnd! Out 5 nmos_a_CDNS_5887047866573 $T=29160 1720 0 90 $X=25260 $Y=1720
.ENDS
***************************************
.SUBCKT cpoly_n_CDNS_588704786656 1 2
** N=2 EP=2 IP=0 FDC=32
M0 1 2 1 cpoly_n w=4.8e-06 l=2e-06 c=5.7348e-14 as=1.44e-13 ad=1.248e-12 ps=2.4e-06 pd=2.13333e-06 sim_w=4.8e-06 m_per_maxw=1 numb_sub_cont=2 nfing=1 $X=620 $Y=200 $D=22
M1 1 2 1 cpoly_n w=4.8e-06 l=2e-06 c=5.7348e-14 as=1.8e-13 ad=1.248e-12 ps=2.4e-06 pd=2.13333e-06 sim_w=4.8e-06 m_per_maxw=1 numb_sub_cont=2 nfing=1 $X=3140 $Y=200 $D=22
M2 1 2 1 cpoly_n w=4.8e-06 l=2e-06 c=5.7348e-14 as=1.8e-13 ad=1.248e-12 ps=2.4e-06 pd=2.13333e-06 sim_w=4.8e-06 m_per_maxw=1 numb_sub_cont=2 nfing=1 $X=5660 $Y=200 $D=22
M3 1 2 1 cpoly_n w=4.8e-06 l=2e-06 c=5.7348e-14 as=1.8e-13 ad=1.248e-12 ps=2.4e-06 pd=2.13333e-06 sim_w=4.8e-06 m_per_maxw=1 numb_sub_cont=2 nfing=1 $X=8180 $Y=200 $D=22
M4 1 2 1 cpoly_n w=4.8e-06 l=2e-06 c=5.7348e-14 as=1.8e-13 ad=1.248e-12 ps=2.4e-06 pd=2.13333e-06 sim_w=4.8e-06 m_per_maxw=1 numb_sub_cont=2 nfing=1 $X=10700 $Y=200 $D=22
M5 1 2 1 cpoly_n w=4.8e-06 l=2e-06 c=5.7348e-14 as=1.8e-13 ad=1.248e-12 ps=2.4e-06 pd=2.13333e-06 sim_w=4.8e-06 m_per_maxw=1 numb_sub_cont=2 nfing=1 $X=13220 $Y=200 $D=22
M6 1 2 1 cpoly_n w=4.8e-06 l=2e-06 c=5.7348e-14 as=1.8e-13 ad=1.248e-12 ps=2.4e-06 pd=2.13333e-06 sim_w=4.8e-06 m_per_maxw=1 numb_sub_cont=2 nfing=1 $X=15740 $Y=200 $D=22
M7 1 2 1 cpoly_n w=4.8e-06 l=2e-06 c=5.7348e-14 as=1.8e-13 ad=1.248e-12 ps=2.4e-06 pd=2.13333e-06 sim_w=4.8e-06 m_per_maxw=1 numb_sub_cont=2 nfing=1 $X=18260 $Y=200 $D=22
M8 1 2 1 cpoly_n w=4.8e-06 l=2e-06 c=5.7348e-14 as=1.8e-13 ad=1.248e-12 ps=2.4e-06 pd=2.13333e-06 sim_w=4.8e-06 m_per_maxw=1 numb_sub_cont=2 nfing=1 $X=20780 $Y=200 $D=22
M9 1 2 1 cpoly_n w=4.8e-06 l=2e-06 c=5.7348e-14 as=1.8e-13 ad=1.248e-12 ps=2.4e-06 pd=2.13333e-06 sim_w=4.8e-06 m_per_maxw=1 numb_sub_cont=2 nfing=1 $X=23300 $Y=200 $D=22
M10 1 2 1 cpoly_n w=4.8e-06 l=2e-06 c=5.7348e-14 as=1.8e-13 ad=1.248e-12 ps=2.4e-06 pd=2.13333e-06 sim_w=4.8e-06 m_per_maxw=1 numb_sub_cont=2 nfing=1 $X=25820 $Y=200 $D=22
M11 1 2 1 cpoly_n w=4.8e-06 l=2e-06 c=5.7348e-14 as=1.8e-13 ad=1.248e-12 ps=2.4e-06 pd=2.13333e-06 sim_w=4.8e-06 m_per_maxw=1 numb_sub_cont=2 nfing=1 $X=28340 $Y=200 $D=22
M12 1 2 1 cpoly_n w=4.8e-06 l=2e-06 c=5.7348e-14 as=1.8e-13 ad=1.248e-12 ps=2.4e-06 pd=2.13333e-06 sim_w=4.8e-06 m_per_maxw=1 numb_sub_cont=2 nfing=1 $X=30860 $Y=200 $D=22
M13 1 2 1 cpoly_n w=4.8e-06 l=2e-06 c=5.7348e-14 as=1.8e-13 ad=1.248e-12 ps=2.4e-06 pd=2.13333e-06 sim_w=4.8e-06 m_per_maxw=1 numb_sub_cont=2 nfing=1 $X=33380 $Y=200 $D=22
M14 1 2 1 cpoly_n w=4.8e-06 l=2e-06 c=5.7348e-14 as=1.8e-13 ad=1.248e-12 ps=2.4e-06 pd=2.13333e-06 sim_w=4.8e-06 m_per_maxw=1 numb_sub_cont=2 nfing=1 $X=35900 $Y=200 $D=22
M15 1 2 1 cpoly_n w=4.8e-06 l=2e-06 c=5.7348e-14 as=1.8e-13 ad=1.248e-12 ps=2.4e-06 pd=2.13333e-06 sim_w=4.8e-06 m_per_maxw=1 numb_sub_cont=2 nfing=1 $X=38420 $Y=200 $D=22
M16 1 2 1 cpoly_n w=4.8e-06 l=2e-06 c=5.7348e-14 as=1.8e-13 ad=1.248e-12 ps=2.4e-06 pd=2.13333e-06 sim_w=4.8e-06 m_per_maxw=1 numb_sub_cont=2 nfing=1 $X=40940 $Y=200 $D=22
M17 1 2 1 cpoly_n w=4.8e-06 l=2e-06 c=5.7348e-14 as=1.8e-13 ad=1.248e-12 ps=2.4e-06 pd=2.13333e-06 sim_w=4.8e-06 m_per_maxw=1 numb_sub_cont=2 nfing=1 $X=43460 $Y=200 $D=22
M18 1 2 1 cpoly_n w=4.8e-06 l=2e-06 c=5.7348e-14 as=1.8e-13 ad=1.248e-12 ps=2.4e-06 pd=2.13333e-06 sim_w=4.8e-06 m_per_maxw=1 numb_sub_cont=2 nfing=1 $X=45980 $Y=200 $D=22
M19 1 2 1 cpoly_n w=4.8e-06 l=2e-06 c=5.7348e-14 as=1.8e-13 ad=1.248e-12 ps=2.4e-06 pd=2.13333e-06 sim_w=4.8e-06 m_per_maxw=1 numb_sub_cont=2 nfing=1 $X=48500 $Y=200 $D=22
M20 1 2 1 cpoly_n w=4.8e-06 l=2e-06 c=5.7348e-14 as=1.8e-13 ad=1.248e-12 ps=2.4e-06 pd=2.13333e-06 sim_w=4.8e-06 m_per_maxw=1 numb_sub_cont=2 nfing=1 $X=51020 $Y=200 $D=22
M21 1 2 1 cpoly_n w=4.8e-06 l=2e-06 c=5.7348e-14 as=1.8e-13 ad=1.248e-12 ps=2.4e-06 pd=2.13333e-06 sim_w=4.8e-06 m_per_maxw=1 numb_sub_cont=2 nfing=1 $X=53540 $Y=200 $D=22
M22 1 2 1 cpoly_n w=4.8e-06 l=2e-06 c=5.7348e-14 as=1.8e-13 ad=1.248e-12 ps=2.4e-06 pd=2.13333e-06 sim_w=4.8e-06 m_per_maxw=1 numb_sub_cont=2 nfing=1 $X=56060 $Y=200 $D=22
M23 1 2 1 cpoly_n w=4.8e-06 l=2e-06 c=5.7348e-14 as=1.8e-13 ad=1.248e-12 ps=2.4e-06 pd=2.13333e-06 sim_w=4.8e-06 m_per_maxw=1 numb_sub_cont=2 nfing=1 $X=58580 $Y=200 $D=22
M24 1 2 1 cpoly_n w=4.8e-06 l=2e-06 c=5.7348e-14 as=1.8e-13 ad=1.248e-12 ps=2.4e-06 pd=2.13333e-06 sim_w=4.8e-06 m_per_maxw=1 numb_sub_cont=2 nfing=1 $X=61100 $Y=200 $D=22
M25 1 2 1 cpoly_n w=4.8e-06 l=2e-06 c=5.7348e-14 as=1.8e-13 ad=1.248e-12 ps=2.4e-06 pd=2.13333e-06 sim_w=4.8e-06 m_per_maxw=1 numb_sub_cont=2 nfing=1 $X=63620 $Y=200 $D=22
M26 1 2 1 cpoly_n w=4.8e-06 l=2e-06 c=5.7348e-14 as=1.8e-13 ad=1.248e-12 ps=2.4e-06 pd=2.13333e-06 sim_w=4.8e-06 m_per_maxw=1 numb_sub_cont=2 nfing=1 $X=66140 $Y=200 $D=22
M27 1 2 1 cpoly_n w=4.8e-06 l=2e-06 c=5.7348e-14 as=1.8e-13 ad=1.248e-12 ps=2.4e-06 pd=2.13333e-06 sim_w=4.8e-06 m_per_maxw=1 numb_sub_cont=2 nfing=1 $X=68660 $Y=200 $D=22
M28 1 2 1 cpoly_n w=4.8e-06 l=2e-06 c=5.7348e-14 as=1.8e-13 ad=1.248e-12 ps=2.4e-06 pd=2.13333e-06 sim_w=4.8e-06 m_per_maxw=1 numb_sub_cont=2 nfing=1 $X=71180 $Y=200 $D=22
M29 1 2 1 cpoly_n w=4.8e-06 l=2e-06 c=5.7348e-14 as=1.8e-13 ad=1.248e-12 ps=2.4e-06 pd=2.13333e-06 sim_w=4.8e-06 m_per_maxw=1 numb_sub_cont=2 nfing=1 $X=73700 $Y=200 $D=22
M30 1 2 1 cpoly_n w=4.8e-06 l=2e-06 c=5.7348e-14 as=1.8e-13 ad=1.248e-12 ps=2.4e-06 pd=2.13333e-06 sim_w=4.8e-06 m_per_maxw=1 numb_sub_cont=2 nfing=1 $X=76220 $Y=200 $D=22
M31 1 2 1 cpoly_n w=4.8e-06 l=2e-06 c=5.7348e-14 as=1.44e-13 ad=1.248e-12 ps=2.4e-06 pd=2.13333e-06 sim_w=4.8e-06 m_per_maxw=1 numb_sub_cont=2 nfing=1 $X=78740 $Y=200 $D=22
.ENDS
***************************************
.SUBCKT cpoly_p_CDNS_588704786655 1 2
** N=2 EP=2 IP=0 FDC=32
M0 1 2 1 cpoly_p w=4.4e-06 l=2e-06 c=5.841e-14 as=1.584e-13 ad=7.488e-13 ps=1.44e-06 pd=1.152e-06 sim_w=2.88e-06 m_per_maxw=1.52778 numb_sub_cont=3 nfing=1 $X=620 $Y=200 $D=21
M1 1 2 1 cpoly_p w=4.4e-06 l=2e-06 c=5.841e-14 as=2.016e-13 ad=7.488e-13 ps=1.44e-06 pd=1.152e-06 sim_w=2.88e-06 m_per_maxw=1.52778 numb_sub_cont=3 nfing=1 $X=3140 $Y=200 $D=21
M2 1 2 1 cpoly_p w=4.4e-06 l=2e-06 c=5.841e-14 as=2.016e-13 ad=7.488e-13 ps=1.44e-06 pd=1.152e-06 sim_w=2.88e-06 m_per_maxw=1.52778 numb_sub_cont=3 nfing=1 $X=5660 $Y=200 $D=21
M3 1 2 1 cpoly_p w=4.4e-06 l=2e-06 c=5.841e-14 as=2.016e-13 ad=7.488e-13 ps=1.44e-06 pd=1.152e-06 sim_w=2.88e-06 m_per_maxw=1.52778 numb_sub_cont=3 nfing=1 $X=8180 $Y=200 $D=21
M4 1 2 1 cpoly_p w=4.4e-06 l=2e-06 c=5.841e-14 as=2.016e-13 ad=7.488e-13 ps=1.44e-06 pd=1.152e-06 sim_w=2.88e-06 m_per_maxw=1.52778 numb_sub_cont=3 nfing=1 $X=10700 $Y=200 $D=21
M5 1 2 1 cpoly_p w=4.4e-06 l=2e-06 c=5.841e-14 as=2.016e-13 ad=7.488e-13 ps=1.44e-06 pd=1.152e-06 sim_w=2.88e-06 m_per_maxw=1.52778 numb_sub_cont=3 nfing=1 $X=13220 $Y=200 $D=21
M6 1 2 1 cpoly_p w=4.4e-06 l=2e-06 c=5.841e-14 as=2.016e-13 ad=7.488e-13 ps=1.44e-06 pd=1.152e-06 sim_w=2.88e-06 m_per_maxw=1.52778 numb_sub_cont=3 nfing=1 $X=15740 $Y=200 $D=21
M7 1 2 1 cpoly_p w=4.4e-06 l=2e-06 c=5.841e-14 as=2.016e-13 ad=7.488e-13 ps=1.44e-06 pd=1.152e-06 sim_w=2.88e-06 m_per_maxw=1.52778 numb_sub_cont=3 nfing=1 $X=18260 $Y=200 $D=21
M8 1 2 1 cpoly_p w=4.4e-06 l=2e-06 c=5.841e-14 as=2.016e-13 ad=7.488e-13 ps=1.44e-06 pd=1.152e-06 sim_w=2.88e-06 m_per_maxw=1.52778 numb_sub_cont=3 nfing=1 $X=20780 $Y=200 $D=21
M9 1 2 1 cpoly_p w=4.4e-06 l=2e-06 c=5.841e-14 as=2.016e-13 ad=7.488e-13 ps=1.44e-06 pd=1.152e-06 sim_w=2.88e-06 m_per_maxw=1.52778 numb_sub_cont=3 nfing=1 $X=23300 $Y=200 $D=21
M10 1 2 1 cpoly_p w=4.4e-06 l=2e-06 c=5.841e-14 as=2.016e-13 ad=7.488e-13 ps=1.44e-06 pd=1.152e-06 sim_w=2.88e-06 m_per_maxw=1.52778 numb_sub_cont=3 nfing=1 $X=25820 $Y=200 $D=21
M11 1 2 1 cpoly_p w=4.4e-06 l=2e-06 c=5.841e-14 as=2.016e-13 ad=7.488e-13 ps=1.44e-06 pd=1.152e-06 sim_w=2.88e-06 m_per_maxw=1.52778 numb_sub_cont=3 nfing=1 $X=28340 $Y=200 $D=21
M12 1 2 1 cpoly_p w=4.4e-06 l=2e-06 c=5.841e-14 as=2.016e-13 ad=7.488e-13 ps=1.44e-06 pd=1.152e-06 sim_w=2.88e-06 m_per_maxw=1.52778 numb_sub_cont=3 nfing=1 $X=30860 $Y=200 $D=21
M13 1 2 1 cpoly_p w=4.4e-06 l=2e-06 c=5.841e-14 as=2.016e-13 ad=7.488e-13 ps=1.44e-06 pd=1.152e-06 sim_w=2.88e-06 m_per_maxw=1.52778 numb_sub_cont=3 nfing=1 $X=33380 $Y=200 $D=21
M14 1 2 1 cpoly_p w=4.4e-06 l=2e-06 c=5.841e-14 as=2.016e-13 ad=7.488e-13 ps=1.44e-06 pd=1.152e-06 sim_w=2.88e-06 m_per_maxw=1.52778 numb_sub_cont=3 nfing=1 $X=35900 $Y=200 $D=21
M15 1 2 1 cpoly_p w=4.4e-06 l=2e-06 c=5.841e-14 as=2.016e-13 ad=7.488e-13 ps=1.44e-06 pd=1.152e-06 sim_w=2.88e-06 m_per_maxw=1.52778 numb_sub_cont=3 nfing=1 $X=38420 $Y=200 $D=21
M16 1 2 1 cpoly_p w=4.4e-06 l=2e-06 c=5.841e-14 as=2.016e-13 ad=7.488e-13 ps=1.44e-06 pd=1.152e-06 sim_w=2.88e-06 m_per_maxw=1.52778 numb_sub_cont=3 nfing=1 $X=40940 $Y=200 $D=21
M17 1 2 1 cpoly_p w=4.4e-06 l=2e-06 c=5.841e-14 as=2.016e-13 ad=7.488e-13 ps=1.44e-06 pd=1.152e-06 sim_w=2.88e-06 m_per_maxw=1.52778 numb_sub_cont=3 nfing=1 $X=43460 $Y=200 $D=21
M18 1 2 1 cpoly_p w=4.4e-06 l=2e-06 c=5.841e-14 as=2.016e-13 ad=7.488e-13 ps=1.44e-06 pd=1.152e-06 sim_w=2.88e-06 m_per_maxw=1.52778 numb_sub_cont=3 nfing=1 $X=45980 $Y=200 $D=21
M19 1 2 1 cpoly_p w=4.4e-06 l=2e-06 c=5.841e-14 as=2.016e-13 ad=7.488e-13 ps=1.44e-06 pd=1.152e-06 sim_w=2.88e-06 m_per_maxw=1.52778 numb_sub_cont=3 nfing=1 $X=48500 $Y=200 $D=21
M20 1 2 1 cpoly_p w=4.4e-06 l=2e-06 c=5.841e-14 as=2.016e-13 ad=7.488e-13 ps=1.44e-06 pd=1.152e-06 sim_w=2.88e-06 m_per_maxw=1.52778 numb_sub_cont=3 nfing=1 $X=51020 $Y=200 $D=21
M21 1 2 1 cpoly_p w=4.4e-06 l=2e-06 c=5.841e-14 as=2.016e-13 ad=7.488e-13 ps=1.44e-06 pd=1.152e-06 sim_w=2.88e-06 m_per_maxw=1.52778 numb_sub_cont=3 nfing=1 $X=53540 $Y=200 $D=21
M22 1 2 1 cpoly_p w=4.4e-06 l=2e-06 c=5.841e-14 as=2.016e-13 ad=7.488e-13 ps=1.44e-06 pd=1.152e-06 sim_w=2.88e-06 m_per_maxw=1.52778 numb_sub_cont=3 nfing=1 $X=56060 $Y=200 $D=21
M23 1 2 1 cpoly_p w=4.4e-06 l=2e-06 c=5.841e-14 as=2.016e-13 ad=7.488e-13 ps=1.44e-06 pd=1.152e-06 sim_w=2.88e-06 m_per_maxw=1.52778 numb_sub_cont=3 nfing=1 $X=58580 $Y=200 $D=21
M24 1 2 1 cpoly_p w=4.4e-06 l=2e-06 c=5.841e-14 as=2.016e-13 ad=7.488e-13 ps=1.44e-06 pd=1.152e-06 sim_w=2.88e-06 m_per_maxw=1.52778 numb_sub_cont=3 nfing=1 $X=61100 $Y=200 $D=21
M25 1 2 1 cpoly_p w=4.4e-06 l=2e-06 c=5.841e-14 as=2.016e-13 ad=7.488e-13 ps=1.44e-06 pd=1.152e-06 sim_w=2.88e-06 m_per_maxw=1.52778 numb_sub_cont=3 nfing=1 $X=63620 $Y=200 $D=21
M26 1 2 1 cpoly_p w=4.4e-06 l=2e-06 c=5.841e-14 as=2.016e-13 ad=7.488e-13 ps=1.44e-06 pd=1.152e-06 sim_w=2.88e-06 m_per_maxw=1.52778 numb_sub_cont=3 nfing=1 $X=66140 $Y=200 $D=21
M27 1 2 1 cpoly_p w=4.4e-06 l=2e-06 c=5.841e-14 as=2.016e-13 ad=7.488e-13 ps=1.44e-06 pd=1.152e-06 sim_w=2.88e-06 m_per_maxw=1.52778 numb_sub_cont=3 nfing=1 $X=68660 $Y=200 $D=21
M28 1 2 1 cpoly_p w=4.4e-06 l=2e-06 c=5.841e-14 as=2.016e-13 ad=7.488e-13 ps=1.44e-06 pd=1.152e-06 sim_w=2.88e-06 m_per_maxw=1.52778 numb_sub_cont=3 nfing=1 $X=71180 $Y=200 $D=21
M29 1 2 1 cpoly_p w=4.4e-06 l=2e-06 c=5.841e-14 as=2.016e-13 ad=7.488e-13 ps=1.44e-06 pd=1.152e-06 sim_w=2.88e-06 m_per_maxw=1.52778 numb_sub_cont=3 nfing=1 $X=73700 $Y=200 $D=21
M30 1 2 1 cpoly_p w=4.4e-06 l=2e-06 c=5.841e-14 as=2.016e-13 ad=7.488e-13 ps=1.44e-06 pd=1.152e-06 sim_w=2.88e-06 m_per_maxw=1.52778 numb_sub_cont=3 nfing=1 $X=76220 $Y=200 $D=21
M31 1 2 1 cpoly_p w=4.4e-06 l=2e-06 c=5.841e-14 as=1.584e-13 ad=7.488e-13 ps=1.44e-06 pd=1.152e-06 sim_w=2.88e-06 m_per_maxw=1.52778 numb_sub_cont=3 nfing=1 $X=78740 $Y=200 $D=21
.ENDS
***************************************
.SUBCKT cpoly_p_CDNS_588704786653 1 2
** N=2 EP=2 IP=0 FDC=32
M0 1 2 1 cpoly_p w=6e-06 l=2e-06 c=8.0712e-14 as=1.68e-13 ad=7.488e-13 ps=1.44e-06 pd=1.13684e-06 sim_w=2.88e-06 m_per_maxw=2.08333 numb_sub_cont=4 nfing=1 $X=620 $Y=200 $D=21
M1 1 2 1 cpoly_p w=6e-06 l=2e-06 c=8.0712e-14 as=2.1408e-13 ad=7.488e-13 ps=1.44e-06 pd=1.13684e-06 sim_w=2.88e-06 m_per_maxw=2.08333 numb_sub_cont=4 nfing=1 $X=3140 $Y=200 $D=21
M2 1 2 1 cpoly_p w=6e-06 l=2e-06 c=8.0712e-14 as=2.1408e-13 ad=7.488e-13 ps=1.44e-06 pd=1.13684e-06 sim_w=2.88e-06 m_per_maxw=2.08333 numb_sub_cont=4 nfing=1 $X=5660 $Y=200 $D=21
M3 1 2 1 cpoly_p w=6e-06 l=2e-06 c=8.0712e-14 as=2.1408e-13 ad=7.488e-13 ps=1.44e-06 pd=1.13684e-06 sim_w=2.88e-06 m_per_maxw=2.08333 numb_sub_cont=4 nfing=1 $X=8180 $Y=200 $D=21
M4 1 2 1 cpoly_p w=6e-06 l=2e-06 c=8.0712e-14 as=2.1408e-13 ad=7.488e-13 ps=1.44e-06 pd=1.13684e-06 sim_w=2.88e-06 m_per_maxw=2.08333 numb_sub_cont=4 nfing=1 $X=10700 $Y=200 $D=21
M5 1 2 1 cpoly_p w=6e-06 l=2e-06 c=8.0712e-14 as=2.1408e-13 ad=7.488e-13 ps=1.44e-06 pd=1.13684e-06 sim_w=2.88e-06 m_per_maxw=2.08333 numb_sub_cont=4 nfing=1 $X=13220 $Y=200 $D=21
M6 1 2 1 cpoly_p w=6e-06 l=2e-06 c=8.0712e-14 as=2.1408e-13 ad=7.488e-13 ps=1.44e-06 pd=1.13684e-06 sim_w=2.88e-06 m_per_maxw=2.08333 numb_sub_cont=4 nfing=1 $X=15740 $Y=200 $D=21
M7 1 2 1 cpoly_p w=6e-06 l=2e-06 c=8.0712e-14 as=2.1408e-13 ad=7.488e-13 ps=1.44e-06 pd=1.13684e-06 sim_w=2.88e-06 m_per_maxw=2.08333 numb_sub_cont=4 nfing=1 $X=18260 $Y=200 $D=21
M8 1 2 1 cpoly_p w=6e-06 l=2e-06 c=8.0712e-14 as=2.1408e-13 ad=7.488e-13 ps=1.44e-06 pd=1.13684e-06 sim_w=2.88e-06 m_per_maxw=2.08333 numb_sub_cont=4 nfing=1 $X=20780 $Y=200 $D=21
M9 1 2 1 cpoly_p w=6e-06 l=2e-06 c=8.0712e-14 as=2.1408e-13 ad=7.488e-13 ps=1.44e-06 pd=1.13684e-06 sim_w=2.88e-06 m_per_maxw=2.08333 numb_sub_cont=4 nfing=1 $X=23300 $Y=200 $D=21
M10 1 2 1 cpoly_p w=6e-06 l=2e-06 c=8.0712e-14 as=2.1408e-13 ad=7.488e-13 ps=1.44e-06 pd=1.13684e-06 sim_w=2.88e-06 m_per_maxw=2.08333 numb_sub_cont=4 nfing=1 $X=25820 $Y=200 $D=21
M11 1 2 1 cpoly_p w=6e-06 l=2e-06 c=8.0712e-14 as=2.1408e-13 ad=7.488e-13 ps=1.44e-06 pd=1.13684e-06 sim_w=2.88e-06 m_per_maxw=2.08333 numb_sub_cont=4 nfing=1 $X=28340 $Y=200 $D=21
M12 1 2 1 cpoly_p w=6e-06 l=2e-06 c=8.0712e-14 as=2.1408e-13 ad=7.488e-13 ps=1.44e-06 pd=1.13684e-06 sim_w=2.88e-06 m_per_maxw=2.08333 numb_sub_cont=4 nfing=1 $X=30860 $Y=200 $D=21
M13 1 2 1 cpoly_p w=6e-06 l=2e-06 c=8.0712e-14 as=2.1408e-13 ad=7.488e-13 ps=1.44e-06 pd=1.13684e-06 sim_w=2.88e-06 m_per_maxw=2.08333 numb_sub_cont=4 nfing=1 $X=33380 $Y=200 $D=21
M14 1 2 1 cpoly_p w=6e-06 l=2e-06 c=8.0712e-14 as=2.1408e-13 ad=7.488e-13 ps=1.44e-06 pd=1.13684e-06 sim_w=2.88e-06 m_per_maxw=2.08333 numb_sub_cont=4 nfing=1 $X=35900 $Y=200 $D=21
M15 1 2 1 cpoly_p w=6e-06 l=2e-06 c=8.0712e-14 as=2.1408e-13 ad=7.488e-13 ps=1.44e-06 pd=1.13684e-06 sim_w=2.88e-06 m_per_maxw=2.08333 numb_sub_cont=4 nfing=1 $X=38420 $Y=200 $D=21
M16 1 2 1 cpoly_p w=6e-06 l=2e-06 c=8.0712e-14 as=2.1408e-13 ad=7.488e-13 ps=1.44e-06 pd=1.13684e-06 sim_w=2.88e-06 m_per_maxw=2.08333 numb_sub_cont=4 nfing=1 $X=40940 $Y=200 $D=21
M17 1 2 1 cpoly_p w=6e-06 l=2e-06 c=8.0712e-14 as=2.1408e-13 ad=7.488e-13 ps=1.44e-06 pd=1.13684e-06 sim_w=2.88e-06 m_per_maxw=2.08333 numb_sub_cont=4 nfing=1 $X=43460 $Y=200 $D=21
M18 1 2 1 cpoly_p w=6e-06 l=2e-06 c=8.0712e-14 as=2.1408e-13 ad=7.488e-13 ps=1.44e-06 pd=1.13684e-06 sim_w=2.88e-06 m_per_maxw=2.08333 numb_sub_cont=4 nfing=1 $X=45980 $Y=200 $D=21
M19 1 2 1 cpoly_p w=6e-06 l=2e-06 c=8.0712e-14 as=2.1408e-13 ad=7.488e-13 ps=1.44e-06 pd=1.13684e-06 sim_w=2.88e-06 m_per_maxw=2.08333 numb_sub_cont=4 nfing=1 $X=48500 $Y=200 $D=21
M20 1 2 1 cpoly_p w=6e-06 l=2e-06 c=8.0712e-14 as=2.1408e-13 ad=7.488e-13 ps=1.44e-06 pd=1.13684e-06 sim_w=2.88e-06 m_per_maxw=2.08333 numb_sub_cont=4 nfing=1 $X=51020 $Y=200 $D=21
M21 1 2 1 cpoly_p w=6e-06 l=2e-06 c=8.0712e-14 as=2.1408e-13 ad=7.488e-13 ps=1.44e-06 pd=1.13684e-06 sim_w=2.88e-06 m_per_maxw=2.08333 numb_sub_cont=4 nfing=1 $X=53540 $Y=200 $D=21
M22 1 2 1 cpoly_p w=6e-06 l=2e-06 c=8.0712e-14 as=2.1408e-13 ad=7.488e-13 ps=1.44e-06 pd=1.13684e-06 sim_w=2.88e-06 m_per_maxw=2.08333 numb_sub_cont=4 nfing=1 $X=56060 $Y=200 $D=21
M23 1 2 1 cpoly_p w=6e-06 l=2e-06 c=8.0712e-14 as=2.1408e-13 ad=7.488e-13 ps=1.44e-06 pd=1.13684e-06 sim_w=2.88e-06 m_per_maxw=2.08333 numb_sub_cont=4 nfing=1 $X=58580 $Y=200 $D=21
M24 1 2 1 cpoly_p w=6e-06 l=2e-06 c=8.0712e-14 as=2.1408e-13 ad=7.488e-13 ps=1.44e-06 pd=1.13684e-06 sim_w=2.88e-06 m_per_maxw=2.08333 numb_sub_cont=4 nfing=1 $X=61100 $Y=200 $D=21
M25 1 2 1 cpoly_p w=6e-06 l=2e-06 c=8.0712e-14 as=2.1408e-13 ad=7.488e-13 ps=1.44e-06 pd=1.13684e-06 sim_w=2.88e-06 m_per_maxw=2.08333 numb_sub_cont=4 nfing=1 $X=63620 $Y=200 $D=21
M26 1 2 1 cpoly_p w=6e-06 l=2e-06 c=8.0712e-14 as=2.1408e-13 ad=7.488e-13 ps=1.44e-06 pd=1.13684e-06 sim_w=2.88e-06 m_per_maxw=2.08333 numb_sub_cont=4 nfing=1 $X=66140 $Y=200 $D=21
M27 1 2 1 cpoly_p w=6e-06 l=2e-06 c=8.0712e-14 as=2.1408e-13 ad=7.488e-13 ps=1.44e-06 pd=1.13684e-06 sim_w=2.88e-06 m_per_maxw=2.08333 numb_sub_cont=4 nfing=1 $X=68660 $Y=200 $D=21
M28 1 2 1 cpoly_p w=6e-06 l=2e-06 c=8.0712e-14 as=2.1408e-13 ad=7.488e-13 ps=1.44e-06 pd=1.13684e-06 sim_w=2.88e-06 m_per_maxw=2.08333 numb_sub_cont=4 nfing=1 $X=71180 $Y=200 $D=21
M29 1 2 1 cpoly_p w=6e-06 l=2e-06 c=8.0712e-14 as=2.1408e-13 ad=7.488e-13 ps=1.44e-06 pd=1.13684e-06 sim_w=2.88e-06 m_per_maxw=2.08333 numb_sub_cont=4 nfing=1 $X=73700 $Y=200 $D=21
M30 1 2 1 cpoly_p w=6e-06 l=2e-06 c=8.0712e-14 as=2.1408e-13 ad=7.488e-13 ps=1.44e-06 pd=1.13684e-06 sim_w=2.88e-06 m_per_maxw=2.08333 numb_sub_cont=4 nfing=1 $X=76220 $Y=200 $D=21
M31 1 2 1 cpoly_p w=6e-06 l=2e-06 c=8.0712e-14 as=1.68e-13 ad=7.488e-13 ps=1.44e-06 pd=1.13684e-06 sim_w=2.88e-06 m_per_maxw=2.08333 numb_sub_cont=4 nfing=1 $X=78740 $Y=200 $D=21
.ENDS
***************************************
.SUBCKT Fill_Dec_X512 vdd! gnd!
** N=2 EP=2 IP=10 FDC=192
M0 vdd! gnd! vdd! cpoly_n w=6e-06 l=2e-06 c=7.5402e-14 as=2.4e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.4338e-06 sim_w=5.76e-06 m_per_maxw=1.04167 numb_sub_cont=3 nfing=1 $X=1360 $Y=47080 $D=22
M1 vdd! gnd! vdd! cpoly_n w=6e-06 l=2e-06 c=7.5402e-14 as=3.0336e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.4338e-06 sim_w=5.76e-06 m_per_maxw=1.04167 numb_sub_cont=3 nfing=1 $X=3880 $Y=47080 $D=22
M2 vdd! gnd! vdd! cpoly_n w=6e-06 l=2e-06 c=7.5402e-14 as=3.0336e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.4338e-06 sim_w=5.76e-06 m_per_maxw=1.04167 numb_sub_cont=3 nfing=1 $X=6400 $Y=47080 $D=22
M3 vdd! gnd! vdd! cpoly_n w=6e-06 l=2e-06 c=7.5402e-14 as=3.0336e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.4338e-06 sim_w=5.76e-06 m_per_maxw=1.04167 numb_sub_cont=3 nfing=1 $X=8920 $Y=47080 $D=22
M4 vdd! gnd! vdd! cpoly_n w=6e-06 l=2e-06 c=7.5402e-14 as=3.0336e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.4338e-06 sim_w=5.76e-06 m_per_maxw=1.04167 numb_sub_cont=3 nfing=1 $X=11440 $Y=47080 $D=22
M5 vdd! gnd! vdd! cpoly_n w=6e-06 l=2e-06 c=7.5402e-14 as=3.0336e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.4338e-06 sim_w=5.76e-06 m_per_maxw=1.04167 numb_sub_cont=3 nfing=1 $X=13960 $Y=47080 $D=22
M6 vdd! gnd! vdd! cpoly_n w=6e-06 l=2e-06 c=7.5402e-14 as=3.0336e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.4338e-06 sim_w=5.76e-06 m_per_maxw=1.04167 numb_sub_cont=3 nfing=1 $X=16480 $Y=47080 $D=22
M7 vdd! gnd! vdd! cpoly_n w=6e-06 l=2e-06 c=7.5402e-14 as=3.0336e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.4338e-06 sim_w=5.76e-06 m_per_maxw=1.04167 numb_sub_cont=3 nfing=1 $X=19000 $Y=47080 $D=22
M8 vdd! gnd! vdd! cpoly_n w=6e-06 l=2e-06 c=7.5402e-14 as=3.0336e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.4338e-06 sim_w=5.76e-06 m_per_maxw=1.04167 numb_sub_cont=3 nfing=1 $X=21520 $Y=47080 $D=22
M9 vdd! gnd! vdd! cpoly_n w=6e-06 l=2e-06 c=7.5402e-14 as=3.0336e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.4338e-06 sim_w=5.76e-06 m_per_maxw=1.04167 numb_sub_cont=3 nfing=1 $X=24040 $Y=47080 $D=22
M10 vdd! gnd! vdd! cpoly_n w=6e-06 l=2e-06 c=7.5402e-14 as=3.0336e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.4338e-06 sim_w=5.76e-06 m_per_maxw=1.04167 numb_sub_cont=3 nfing=1 $X=26560 $Y=47080 $D=22
M11 vdd! gnd! vdd! cpoly_n w=6e-06 l=2e-06 c=7.5402e-14 as=3.0336e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.4338e-06 sim_w=5.76e-06 m_per_maxw=1.04167 numb_sub_cont=3 nfing=1 $X=29080 $Y=47080 $D=22
M12 vdd! gnd! vdd! cpoly_n w=6e-06 l=2e-06 c=7.5402e-14 as=3.0336e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.4338e-06 sim_w=5.76e-06 m_per_maxw=1.04167 numb_sub_cont=3 nfing=1 $X=31600 $Y=47080 $D=22
M13 vdd! gnd! vdd! cpoly_n w=6e-06 l=2e-06 c=7.5402e-14 as=3.0336e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.4338e-06 sim_w=5.76e-06 m_per_maxw=1.04167 numb_sub_cont=3 nfing=1 $X=34120 $Y=47080 $D=22
M14 vdd! gnd! vdd! cpoly_n w=6e-06 l=2e-06 c=7.5402e-14 as=3.0336e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.4338e-06 sim_w=5.76e-06 m_per_maxw=1.04167 numb_sub_cont=3 nfing=1 $X=36640 $Y=47080 $D=22
M15 vdd! gnd! vdd! cpoly_n w=6e-06 l=2e-06 c=7.5402e-14 as=3.0336e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.4338e-06 sim_w=5.76e-06 m_per_maxw=1.04167 numb_sub_cont=3 nfing=1 $X=39160 $Y=47080 $D=22
M16 vdd! gnd! vdd! cpoly_n w=6e-06 l=2e-06 c=7.5402e-14 as=3.0336e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.4338e-06 sim_w=5.76e-06 m_per_maxw=1.04167 numb_sub_cont=3 nfing=1 $X=41680 $Y=47080 $D=22
M17 vdd! gnd! vdd! cpoly_n w=6e-06 l=2e-06 c=7.5402e-14 as=3.0336e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.4338e-06 sim_w=5.76e-06 m_per_maxw=1.04167 numb_sub_cont=3 nfing=1 $X=44200 $Y=47080 $D=22
M18 vdd! gnd! vdd! cpoly_n w=6e-06 l=2e-06 c=7.5402e-14 as=3.0336e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.4338e-06 sim_w=5.76e-06 m_per_maxw=1.04167 numb_sub_cont=3 nfing=1 $X=46720 $Y=47080 $D=22
M19 vdd! gnd! vdd! cpoly_n w=6e-06 l=2e-06 c=7.5402e-14 as=3.0336e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.4338e-06 sim_w=5.76e-06 m_per_maxw=1.04167 numb_sub_cont=3 nfing=1 $X=49240 $Y=47080 $D=22
M20 vdd! gnd! vdd! cpoly_n w=6e-06 l=2e-06 c=7.5402e-14 as=3.0336e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.4338e-06 sim_w=5.76e-06 m_per_maxw=1.04167 numb_sub_cont=3 nfing=1 $X=51760 $Y=47080 $D=22
M21 vdd! gnd! vdd! cpoly_n w=6e-06 l=2e-06 c=7.5402e-14 as=3.0336e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.4338e-06 sim_w=5.76e-06 m_per_maxw=1.04167 numb_sub_cont=3 nfing=1 $X=54280 $Y=47080 $D=22
M22 vdd! gnd! vdd! cpoly_n w=6e-06 l=2e-06 c=7.5402e-14 as=3.0336e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.4338e-06 sim_w=5.76e-06 m_per_maxw=1.04167 numb_sub_cont=3 nfing=1 $X=56800 $Y=47080 $D=22
M23 vdd! gnd! vdd! cpoly_n w=6e-06 l=2e-06 c=7.5402e-14 as=3.0336e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.4338e-06 sim_w=5.76e-06 m_per_maxw=1.04167 numb_sub_cont=3 nfing=1 $X=59320 $Y=47080 $D=22
M24 vdd! gnd! vdd! cpoly_n w=6e-06 l=2e-06 c=7.5402e-14 as=3.0336e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.4338e-06 sim_w=5.76e-06 m_per_maxw=1.04167 numb_sub_cont=3 nfing=1 $X=61840 $Y=47080 $D=22
M25 vdd! gnd! vdd! cpoly_n w=6e-06 l=2e-06 c=7.5402e-14 as=3.0336e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.4338e-06 sim_w=5.76e-06 m_per_maxw=1.04167 numb_sub_cont=3 nfing=1 $X=64360 $Y=47080 $D=22
M26 vdd! gnd! vdd! cpoly_n w=6e-06 l=2e-06 c=7.5402e-14 as=3.0336e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.4338e-06 sim_w=5.76e-06 m_per_maxw=1.04167 numb_sub_cont=3 nfing=1 $X=66880 $Y=47080 $D=22
M27 vdd! gnd! vdd! cpoly_n w=6e-06 l=2e-06 c=7.5402e-14 as=3.0336e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.4338e-06 sim_w=5.76e-06 m_per_maxw=1.04167 numb_sub_cont=3 nfing=1 $X=69400 $Y=47080 $D=22
M28 vdd! gnd! vdd! cpoly_n w=6e-06 l=2e-06 c=7.5402e-14 as=3.0336e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.4338e-06 sim_w=5.76e-06 m_per_maxw=1.04167 numb_sub_cont=3 nfing=1 $X=71920 $Y=47080 $D=22
M29 vdd! gnd! vdd! cpoly_n w=6e-06 l=2e-06 c=7.5402e-14 as=3.0336e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.4338e-06 sim_w=5.76e-06 m_per_maxw=1.04167 numb_sub_cont=3 nfing=1 $X=74440 $Y=47080 $D=22
M30 vdd! gnd! vdd! cpoly_n w=6e-06 l=2e-06 c=7.5402e-14 as=3.0336e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.4338e-06 sim_w=5.76e-06 m_per_maxw=1.04167 numb_sub_cont=3 nfing=1 $X=76960 $Y=47080 $D=22
M31 vdd! gnd! vdd! cpoly_n w=6e-06 l=2e-06 c=7.5402e-14 as=2.4e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.4338e-06 sim_w=5.76e-06 m_per_maxw=1.04167 numb_sub_cont=3 nfing=1 $X=79480 $Y=47080 $D=22
X32 vdd! gnd! cpoly_n_CDNS_588704786656 $T=82100 8440 1 180 $X=740 $Y=8440
X33 vdd! gnd! cpoly_n_CDNS_588704786656 $T=82100 27660 1 180 $X=740 $Y=27660
X34 gnd! vdd! cpoly_p_CDNS_588704786655 $T=740 19900 0 0 $X=740 $Y=19900
X35 gnd! vdd! cpoly_p_CDNS_588704786655 $T=740 39120 0 0 $X=740 $Y=39120
X36 gnd! vdd! cpoly_p_CDNS_588704786653 $T=740 56240 0 0 $X=740 $Y=56240
.ENDS
***************************************
.SUBCKT ICV_91 1 2 3
** N=3 EP=3 IP=7 FDC=4
D0 2 1 dn PJ=0.00041 m=1 $X=5220 $Y=0 $D=8
D1 1 3 dn PJ=0.00041 m=1 $X=7720 $Y=0 $D=8
X4 3 1 2 ICV_84 $T=0 0 0 0 $X=-640 $Y=-300
.ENDS
***************************************
.SUBCKT ICV_92 1 2 3
** N=3 EP=3 IP=6 FDC=8
X0 2 3 1 ICV_91 $T=0 0 0 0 $X=-640 $Y=-300
X1 2 3 1 ICV_91 $T=10000 0 0 0 $X=9360 $Y=-300
.ENDS
***************************************
.SUBCKT GND_Core_PAD gnd! GND_PAD vdd!
** N=8 EP=3 IP=21 FDC=115
D0 gnd! vdd! dn PJ=0.00041 m=1 $X=94280 $Y=-99700 $D=9
X1 vdd! gnd! cpoly_n_CDNS_588704786651 $T=520 333340 0 0 $X=520 $Y=333340
X2 gnd! vdd! cpoly_p_CDNS_588704786650 $T=520 320500 0 0 $X=520 $Y=320500
X4 gnd! GND_PAD vdd! ICV_91 $T=84740 -99700 0 0 $X=84100 $Y=-100000
X5 vdd! gnd! GND_PAD ICV_92 $T=4740 -99700 0 0 $X=4100 $Y=-100000
X6 vdd! gnd! GND_PAD ICV_92 $T=24740 -99700 0 0 $X=24100 $Y=-100000
X7 vdd! gnd! GND_PAD ICV_92 $T=44740 -99700 0 0 $X=44100 $Y=-100000
X8 vdd! gnd! GND_PAD ICV_92 $T=64740 -99700 0 0 $X=64100 $Y=-100000
.ENDS
***************************************
.SUBCKT nmos_a_CDNS_5887047866563
** N=2 EP=0 IP=0 FDC=0
*.SEEDPROM
.ENDS
***************************************
.SUBCKT ICV_93 1 2
** N=2 EP=2 IP=4 FDC=2
M0 1 2 1 1 nmos_a L=2e-06 W=9.6e-05 AD=1.2132e-12 AS=2.496e-11 PD=3.033e-06 PS=1.5165e-06 w_cont=5.1e-06 nfing=1 source_num=2 $X=-1900 $Y=200 $D=1
M1 1 2 1 1 nmos_a L=2e-06 W=9.6e-05 AD=1.2132e-12 AS=2.496e-11 PD=3.033e-06 PS=1.5165e-06 w_cont=5.1e-06 nfing=1 source_num=2 $X=620 $Y=200 $D=1
.ENDS
***************************************
.SUBCKT dn_CDNS_5887047866564 1 2
** N=2 EP=2 IP=0 FDC=1
D0 2 1 dn PJ=5e-07 m=1 $X=-460 $Y=0 $D=9
.ENDS
***************************************
.SUBCKT nmos_io_a_CDNS_5887047866565
** N=3 EP=0 IP=0 FDC=0
*.SEEDPROM
.ENDS
***************************************
.SUBCKT nmos_a_CDNS_5887047866562 1 2
** N=2 EP=2 IP=0 FDC=1
M0 1 2 1 1 nmos_a L=2e-06 W=9.4e-05 AD=1.2145e-12 AS=3.76e-11 PD=3.03626e-06 PS=1.51813e-06 w_cont=5.1e-06 nfing=1 source_num=2 $X=620 $Y=200 $D=1
.ENDS
***************************************
.SUBCKT Usub_7V_ESD GND_PAD! Minus3 Minus6_VD 5 UsubVD Minus6 Usub
** N=8 EP=7 IP=48 FDC=25
*.SEEDPROM
M0 Minus6_VD UsubVD Usub Usub nmos_io_a L=2.8e-07 W=7.4e-05 AD=7.12574e-12 AS=2.21449e-13 PD=3.91524e-06 PS=1.95762e-06 w_cont=2.66e-05 nfing=1 $X=620 $Y=200 $D=0
M1 5 Minus6 Minus6_VD Minus6_VD nmos_io_a L=2.8e-07 W=7.4e-05 AD=7.12574e-12 AS=2.21449e-13 PD=3.91524e-06 PS=1.95762e-06 w_cont=2.66e-05 nfing=1 $X=620 $Y=207640 $D=0
M2 5 Minus6 Minus6_VD Minus6_VD nmos_io_a L=2.8e-07 W=7.4e-05 AD=7.12574e-12 AS=2.21449e-13 PD=3.91524e-06 PS=1.95762e-06 w_cont=2.66e-05 nfing=1 $X=620 $Y=311080 $D=0
M3 GND_PAD! Minus3 5 5 nmos_io_a L=2.8e-07 W=7.4e-05 AD=7.12574e-12 AS=2.21449e-13 PD=3.91524e-06 PS=1.95762e-06 w_cont=2.66e-05 nfing=1 $X=6720 $Y=200 $D=0
M4 GND_PAD! Minus3 5 5 nmos_io_a L=2.8e-07 W=7.4e-05 AD=7.12574e-12 AS=2.21449e-13 PD=3.91524e-06 PS=1.95762e-06 w_cont=2.66e-05 nfing=1 $X=6720 $Y=103920 $D=0
M5 GND_PAD! Minus3 5 5 nmos_io_a L=2.8e-07 W=7.4e-05 AD=7.12574e-12 AS=2.21449e-13 PD=3.91524e-06 PS=1.95762e-06 w_cont=2.66e-05 nfing=1 $X=6720 $Y=207640 $D=0
M6 GND_PAD! Minus3 5 5 nmos_io_a L=2.8e-07 W=7.4e-05 AD=7.12574e-12 AS=2.21449e-13 PD=3.91524e-06 PS=1.95762e-06 w_cont=2.66e-05 nfing=1 $X=6720 $Y=311360 $D=0
M7 UsubVD Minus6 UsubVD UsubVD nmos_a L=2e-06 W=9.6e-05 AD=1.2132e-12 AS=3.84e-11 PD=3.033e-06 PS=1.5165e-06 w_cont=5.1e-06 nfing=1 source_num=2 $X=3520 $Y=200 $D=1
D8 Usub UsubVD dn PJ=5e-07 m=1 $X=1780 $Y=101680 $D=9
D9 Minus6_VD Minus6 dn PJ=5e-07 m=1 $X=1780 $Y=205500 $D=9
X11 GND_PAD! Minus3 ICV_93 $T=12200 0 1 180 $X=9000 $Y=0
X12 GND_PAD! Minus3 ICV_93 $T=12200 103720 1 180 $X=9000 $Y=103720
X13 GND_PAD! Minus3 ICV_93 $T=12200 207440 1 180 $X=9000 $Y=207440
X14 GND_PAD! Minus3 ICV_93 $T=12200 311020 1 180 $X=9000 $Y=311020
X15 Minus6 Minus6_VD dn_CDNS_5887047866564 $T=2300 309560 0 180 $X=900 $Y=308760
X16 Minus3 5 dn_CDNS_5887047866564 $T=8400 102180 0 180 $X=7000 $Y=101380
X17 Minus3 5 dn_CDNS_5887047866564 $T=8400 205900 0 180 $X=7000 $Y=205100
X18 Minus3 5 dn_CDNS_5887047866564 $T=8400 309620 0 180 $X=7000 $Y=308820
X27 Minus3 Minus6 nmos_a_CDNS_5887047866562 $T=2900 104300 0 0 $X=2900 $Y=104300
X28 Minus3 Minus6 nmos_a_CDNS_5887047866562 $T=2900 208200 0 0 $X=2900 $Y=208200
X29 Minus3 Minus6 nmos_a_CDNS_5887047866562 $T=2900 311620 0 0 $X=2900 $Y=311620
.ENDS
***************************************
.SUBCKT ICV_94 1 3 4 5 7 8 9
** N=9 EP=7 IP=8 FDC=26
M0 8 4 3 3 nmos_io_a L=2.8e-07 W=7.4e-05 AD=7.12574e-12 AS=2.42621e-13 PD=3.91524e-06 PS=1.95762e-06 w_cont=2.66e-05 nfing=1 $X=620 $Y=103920 $D=0
X1 1 7 8 9 4 5 3 Usub_7V_ESD $T=0 0 0 0 $X=0 $Y=-3160
.ENDS
***************************************
.SUBCKT ICV_95 1 3 4 5 7 8 9
** N=9 EP=7 IP=8 FDC=26
M0 8 4 3 3 nmos_io_a L=2.8e-07 W=7.4e-05 AD=7.12574e-12 AS=2.21449e-13 PD=3.91524e-06 PS=1.95762e-06 w_cont=2.66e-05 nfing=1 $X=620 $Y=103920 $D=0
X1 1 7 8 9 4 5 3 Usub_7V_ESD $T=0 0 0 0 $X=0 $Y=-3160
.ENDS
***************************************
.SUBCKT ICV_96 1 3 4 5 7 8 9
** N=9 EP=7 IP=8 FDC=26
M0 8 4 3 3 nmos_io_a L=2.8e-07 W=7.4e-05 AD=7.12574e-12 AS=2.21449e-13 PD=3.91524e-06 PS=1.95762e-06 w_cont=2.66e-05 nfing=1 $X=620 $Y=103920 $D=0
X1 1 7 8 9 4 5 3 Usub_7V_ESD $T=0 0 0 0 $X=0 $Y=-3160
.ENDS
***************************************
.SUBCKT ICV_97 1 3 4 5 7 8 9
** N=9 EP=7 IP=8 FDC=26
M0 8 4 3 3 nmos_io_a L=2.8e-07 W=7.4e-05 AD=7.12574e-12 AS=2.21449e-13 PD=3.91524e-06 PS=1.95762e-06 w_cont=2.66e-05 nfing=1 $X=620 $Y=103920 $D=0
X1 1 7 8 9 4 5 3 Usub_7V_ESD $T=0 0 0 0 $X=0 $Y=-3160
.ENDS
***************************************
.SUBCKT ICV_98 1 3 4 5 7 8 9
** N=9 EP=7 IP=8 FDC=26
M0 8 4 3 3 nmos_io_a L=2.8e-07 W=7.4e-05 AD=7.12574e-12 AS=2.21449e-13 PD=3.91524e-06 PS=1.95762e-06 w_cont=2.66e-05 nfing=1 $X=620 $Y=103920 $D=0
X1 1 7 8 9 4 5 3 Usub_7V_ESD $T=0 0 0 0 $X=0 $Y=-3160
.ENDS
***************************************
.SUBCKT ICV_99 1 3 4 5 7 8 9
** N=9 EP=7 IP=8 FDC=26
M0 8 4 3 3 nmos_io_a L=2.8e-07 W=7.4e-05 AD=7.12574e-12 AS=2.21449e-13 PD=3.91524e-06 PS=1.95762e-06 w_cont=2.66e-05 nfing=1 $X=620 $Y=103920 $D=0
X1 1 7 8 9 4 5 3 Usub_7V_ESD $T=0 0 0 0 $X=0 $Y=-3160
.ENDS
***************************************
.SUBCKT ICV_100 1 3 4 5 7 8 9
** N=9 EP=7 IP=8 FDC=26
M0 8 4 3 3 nmos_io_a L=2.8e-07 W=7.4e-05 AD=7.12574e-12 AS=2.21449e-13 PD=3.91524e-06 PS=1.95762e-06 w_cont=2.66e-05 nfing=1 $X=620 $Y=103920 $D=0
X1 1 7 8 9 4 5 3 Usub_7V_ESD $T=0 0 0 0 $X=0 $Y=-3160
.ENDS
***************************************
.SUBCKT ICV_101 1 3 4 5 7 8 9
** N=9 EP=7 IP=8 FDC=26
M0 8 4 3 3 nmos_io_a L=2.8e-07 W=7.4e-05 AD=7.12574e-12 AS=2.21449e-13 PD=3.91524e-06 PS=1.95762e-06 w_cont=2.66e-05 nfing=1 $X=620 $Y=103920 $D=0
X1 1 7 8 9 4 5 3 Usub_7V_ESD $T=0 0 0 0 $X=0 $Y=-3160
.ENDS
***************************************
.SUBCKT ICV_102 1 3 4 5 7 8 9
** N=9 EP=7 IP=8 FDC=26
M0 8 4 3 3 nmos_io_a L=2.8e-07 W=7.4e-05 AD=7.12574e-12 AS=2.21449e-13 PD=3.91524e-06 PS=1.95762e-06 w_cont=2.66e-05 nfing=1 $X=620 $Y=103920 $D=0
X1 1 7 8 9 4 5 3 Usub_7V_ESD $T=0 0 0 0 $X=0 $Y=-3160
.ENDS
***************************************
.SUBCKT ICV_103 1 3 4 5 7 8 9
** N=9 EP=7 IP=8 FDC=26
M0 8 4 3 3 nmos_io_a L=2.8e-07 W=7.4e-05 AD=7.12574e-12 AS=2.21449e-13 PD=3.91524e-06 PS=1.95762e-06 w_cont=2.66e-05 nfing=1 $X=620 $Y=103920 $D=0
X1 1 7 8 9 4 5 3 Usub_7V_ESD $T=0 0 0 0 $X=0 $Y=-3160
.ENDS
***************************************
.SUBCKT ICV_104 1 3 4 5 7 8 9
** N=9 EP=7 IP=8 FDC=26
M0 8 4 3 3 nmos_io_a L=2.8e-07 W=7.4e-05 AD=7.12574e-12 AS=2.21449e-13 PD=3.91524e-06 PS=1.95762e-06 w_cont=2.66e-05 nfing=1 $X=620 $Y=103920 $D=0
X1 1 7 8 9 4 5 3 Usub_7V_ESD $T=0 0 0 0 $X=0 $Y=-3160
.ENDS
***************************************
.SUBCKT ICV_105 1 3 4 5 7 8 9
** N=9 EP=7 IP=8 FDC=26
M0 8 4 3 3 nmos_io_a L=2.8e-07 W=7.4e-05 AD=7.12574e-12 AS=2.21449e-13 PD=3.91524e-06 PS=1.95762e-06 w_cont=2.66e-05 nfing=1 $X=620 $Y=103920 $D=0
X1 1 7 8 9 4 5 3 Usub_7V_ESD $T=0 0 0 0 $X=0 $Y=-3160
.ENDS
***************************************
.SUBCKT ICV_106 1 3 4 5 7 8 9
** N=9 EP=7 IP=8 FDC=26
M0 8 4 3 3 nmos_io_a L=2.8e-07 W=7.4e-05 AD=7.12574e-12 AS=2.21449e-13 PD=3.91524e-06 PS=1.95762e-06 w_cont=2.66e-05 nfing=1 $X=620 $Y=103920 $D=0
X1 1 7 8 9 4 5 3 Usub_7V_ESD $T=0 0 0 0 $X=0 $Y=-3160
.ENDS
***************************************
.SUBCKT ICV_107 1 3 4 5 7 8 9
** N=9 EP=7 IP=8 FDC=26
M0 8 4 3 3 nmos_io_a L=2.8e-07 W=7.4e-05 AD=7.12574e-12 AS=2.21449e-13 PD=3.91524e-06 PS=1.95762e-06 w_cont=2.66e-05 nfing=1 $X=620 $Y=103920 $D=0
X1 1 7 8 9 4 5 3 Usub_7V_ESD $T=0 0 0 0 $X=0 $Y=-3160
.ENDS
***************************************
.SUBCKT ICV_108 1 3 4 5 7 8 9
** N=9 EP=7 IP=8 FDC=26
M0 8 4 3 3 nmos_io_a L=2.8e-07 W=7.4e-05 AD=7.12574e-12 AS=2.21449e-13 PD=3.91524e-06 PS=1.95762e-06 w_cont=2.66e-05 nfing=1 $X=620 $Y=103920 $D=0
X1 1 7 8 9 4 5 3 Usub_7V_ESD $T=0 0 0 0 $X=0 $Y=-3160
.ENDS
***************************************
.SUBCKT ICV_109 1 3 4 5 7 8 9
** N=9 EP=7 IP=8 FDC=26
M0 8 4 3 3 nmos_io_a L=2.8e-07 W=7.4e-05 AD=7.12574e-12 AS=2.21449e-13 PD=3.91524e-06 PS=1.95762e-06 w_cont=2.66e-05 nfing=1 $X=620 $Y=103920 $D=0
X1 1 7 8 9 4 5 3 Usub_7V_ESD $T=0 0 0 0 $X=0 $Y=-3160
.ENDS
***************************************
.SUBCKT ICV_110 1 3 4 5 7 8 9
** N=9 EP=7 IP=8 FDC=26
M0 8 4 3 3 nmos_io_a L=2.8e-07 W=7.4e-05 AD=7.12574e-12 AS=2.21449e-13 PD=3.91524e-06 PS=1.95762e-06 w_cont=2.66e-05 nfing=1 $X=620 $Y=103920 $D=0
X1 1 7 8 9 4 5 3 Usub_7V_ESD $T=0 0 0 0 $X=0 $Y=-3160
.ENDS
***************************************
.SUBCKT ICV_111 1 3 4 5 7 8 9
** N=9 EP=7 IP=8 FDC=26
M0 8 4 3 3 nmos_io_a L=2.8e-07 W=7.4e-05 AD=7.12574e-12 AS=2.21449e-13 PD=3.91524e-06 PS=1.95762e-06 w_cont=2.66e-05 nfing=1 $X=620 $Y=103920 $D=0
X1 1 7 8 9 4 5 3 Usub_7V_ESD $T=0 0 0 0 $X=0 $Y=-3160
.ENDS
***************************************
.SUBCKT ICV_112 1 3 4 5 7 8 9
** N=9 EP=7 IP=8 FDC=26
M0 8 4 3 3 nmos_io_a L=2.8e-07 W=7.4e-05 AD=7.12574e-12 AS=2.21449e-13 PD=3.91524e-06 PS=1.95762e-06 w_cont=2.66e-05 nfing=1 $X=620 $Y=103920 $D=0
X1 1 7 8 9 4 5 3 Usub_7V_ESD $T=0 0 0 0 $X=0 $Y=-3160
.ENDS
***************************************
.SUBCKT ICV_113 1 3 4 5 7 8 9
** N=9 EP=7 IP=8 FDC=26
M0 8 4 3 3 nmos_io_a L=2.8e-07 W=7.4e-05 AD=7.12574e-12 AS=2.21449e-13 PD=3.91524e-06 PS=1.95762e-06 w_cont=2.66e-05 nfing=1 $X=620 $Y=103920 $D=0
X1 1 7 8 9 4 5 3 Usub_7V_ESD $T=0 0 0 0 $X=0 $Y=-3160
.ENDS
***************************************
.SUBCKT ICV_114 1 3 4 5 7 8 9
** N=9 EP=7 IP=8 FDC=26
M0 8 4 3 3 nmos_io_a L=2.8e-07 W=7.4e-05 AD=7.12574e-12 AS=2.21449e-13 PD=3.91524e-06 PS=1.95762e-06 w_cont=2.66e-05 nfing=1 $X=620 $Y=103920 $D=0
X1 1 7 8 9 4 5 3 Usub_7V_ESD $T=0 0 0 0 $X=0 $Y=-3160
.ENDS
***************************************
.SUBCKT ICV_115 1 3 4 5 7 8 9
** N=9 EP=7 IP=8 FDC=26
M0 8 4 3 3 nmos_io_a L=2.8e-07 W=7.4e-05 AD=7.12574e-12 AS=2.21449e-13 PD=3.91524e-06 PS=1.95762e-06 w_cont=2.66e-05 nfing=1 $X=620 $Y=103920 $D=0
X1 1 7 8 9 4 5 3 Usub_7V_ESD $T=0 0 0 0 $X=0 $Y=-3160
.ENDS
***************************************
.SUBCKT ICV_116 1 3 4 5 7 8 9
** N=9 EP=7 IP=8 FDC=26
M0 8 4 3 3 nmos_io_a L=2.8e-07 W=7.4e-05 AD=7.12574e-12 AS=2.21449e-13 PD=3.91524e-06 PS=1.95762e-06 w_cont=2.66e-05 nfing=1 $X=620 $Y=103920 $D=0
X1 1 7 8 9 4 5 3 Usub_7V_ESD $T=0 0 0 0 $X=0 $Y=-3160
.ENDS
***************************************
.SUBCKT ICV_117 1 3 4 5 7 8 9
** N=9 EP=7 IP=8 FDC=26
M0 8 4 3 3 nmos_io_a L=2.8e-07 W=7.4e-05 AD=7.12574e-12 AS=2.21449e-13 PD=3.91524e-06 PS=1.95762e-06 w_cont=2.66e-05 nfing=1 $X=620 $Y=103920 $D=0
X1 1 7 8 9 4 5 3 Usub_7V_ESD $T=0 0 0 0 $X=0 $Y=-3160
.ENDS
***************************************
.SUBCKT ICV_118 1 3 4 5 7 8 9
** N=9 EP=7 IP=8 FDC=26
M0 8 4 3 3 nmos_io_a L=2.8e-07 W=7.4e-05 AD=7.12574e-12 AS=2.21449e-13 PD=3.91524e-06 PS=1.95762e-06 w_cont=2.66e-05 nfing=1 $X=620 $Y=103920 $D=0
X1 1 7 8 9 4 5 3 Usub_7V_ESD $T=0 0 0 0 $X=0 $Y=-3160
.ENDS
***************************************
.SUBCKT ICV_119 1 3 4 5 7 8 9
** N=9 EP=7 IP=8 FDC=26
M0 8 4 3 3 nmos_io_a L=2.8e-07 W=7.4e-05 AD=7.12574e-12 AS=2.21449e-13 PD=3.91524e-06 PS=1.95762e-06 w_cont=2.66e-05 nfing=1 $X=620 $Y=103920 $D=0
X1 1 7 8 9 4 5 3 Usub_7V_ESD $T=0 0 0 0 $X=0 $Y=-3160
.ENDS
***************************************
.SUBCKT ICV_120 1 3 4 5 7 8 9
** N=9 EP=7 IP=8 FDC=26
M0 8 4 3 3 nmos_io_a L=2.8e-07 W=7.4e-05 AD=7.12574e-12 AS=2.21449e-13 PD=3.91524e-06 PS=1.95762e-06 w_cont=2.66e-05 nfing=1 $X=620 $Y=103920 $D=0
X1 1 7 8 9 4 5 3 Usub_7V_ESD $T=0 0 0 0 $X=0 $Y=-3160
.ENDS
***************************************
.SUBCKT ICV_121 1 3 4 5 7 8 9
** N=9 EP=7 IP=8 FDC=26
M0 8 4 3 3 nmos_io_a L=2.8e-07 W=7.4e-05 AD=7.12574e-12 AS=2.21449e-13 PD=3.91524e-06 PS=1.95762e-06 w_cont=2.66e-05 nfing=1 $X=620 $Y=103920 $D=0
X1 1 7 8 9 4 5 3 Usub_7V_ESD $T=0 0 0 0 $X=0 $Y=-3160
.ENDS
***************************************
.SUBCKT ICV_122 1 3 4 5 7 8 9
** N=9 EP=7 IP=8 FDC=26
M0 8 4 3 3 nmos_io_a L=2.8e-07 W=7.4e-05 AD=7.12574e-12 AS=2.21449e-13 PD=3.91524e-06 PS=1.95762e-06 w_cont=2.66e-05 nfing=1 $X=620 $Y=103920 $D=0
X1 1 7 8 9 4 5 3 Usub_7V_ESD $T=0 0 0 0 $X=0 $Y=-3160
.ENDS
***************************************
.SUBCKT ICV_123 1 3 4 5 7 8 9
** N=9 EP=7 IP=8 FDC=26
M0 8 4 3 3 nmos_io_a L=2.8e-07 W=7.4e-05 AD=7.12574e-12 AS=2.21449e-13 PD=3.91524e-06 PS=1.95762e-06 w_cont=2.66e-05 nfing=1 $X=620 $Y=103920 $D=0
X1 1 7 8 9 4 5 3 Usub_7V_ESD $T=0 0 0 0 $X=0 $Y=-3160
.ENDS
***************************************
.SUBCKT ICV_124 1 3 4 5 7 8 9
** N=9 EP=7 IP=8 FDC=26
M0 8 4 3 3 nmos_io_a L=2.8e-07 W=7.4e-05 AD=7.12574e-12 AS=2.21449e-13 PD=3.91524e-06 PS=1.95762e-06 w_cont=2.66e-05 nfing=1 $X=620 $Y=103920 $D=0
X1 1 7 8 9 4 5 3 Usub_7V_ESD $T=0 0 0 0 $X=0 $Y=-3160
.ENDS
***************************************
.SUBCKT ICV_125 1 3 4 5 7 8 9
** N=9 EP=7 IP=8 FDC=26
M0 8 4 3 3 nmos_io_a L=2.8e-07 W=7.4e-05 AD=7.12574e-12 AS=2.21449e-13 PD=3.91524e-06 PS=1.95762e-06 w_cont=2.66e-05 nfing=1 $X=620 $Y=103920 $D=0
X1 1 7 8 9 4 5 3 Usub_7V_ESD $T=0 0 0 0 $X=0 $Y=-3160
.ENDS
***************************************
.SUBCKT ICV_126 1 3 4 5 7 8 9
** N=9 EP=7 IP=8 FDC=26
M0 8 4 3 3 nmos_io_a L=2.8e-07 W=7.4e-05 AD=7.12574e-12 AS=2.21449e-13 PD=3.91524e-06 PS=1.95762e-06 w_cont=2.66e-05 nfing=1 $X=620 $Y=103920 $D=0
X1 1 7 8 9 4 5 3 Usub_7V_ESD $T=0 0 0 0 $X=0 $Y=-3160
.ENDS
***************************************
.SUBCKT ICV_127 1 3 4 5 7 8 9
** N=9 EP=7 IP=8 FDC=26
M0 8 4 3 3 nmos_io_a L=2.8e-07 W=7.4e-05 AD=7.12574e-12 AS=2.21449e-13 PD=3.91524e-06 PS=1.95762e-06 w_cont=2.66e-05 nfing=1 $X=620 $Y=103920 $D=0
X1 1 7 8 9 4 5 3 Usub_7V_ESD $T=0 0 0 0 $X=0 $Y=-3160
.ENDS
***************************************
.SUBCKT ICV_128 1 3 4 5 7 8 9
** N=9 EP=7 IP=8 FDC=26
M0 8 4 3 3 nmos_io_a L=2.8e-07 W=7.4e-05 AD=7.12574e-12 AS=2.21449e-13 PD=3.91524e-06 PS=1.95762e-06 w_cont=2.66e-05 nfing=1 $X=620 $Y=103920 $D=0
X1 1 7 8 9 4 5 3 Usub_7V_ESD $T=0 0 0 0 $X=0 $Y=-3160
.ENDS
***************************************
.SUBCKT ICV_129 1 3 4 5 7 8 9
** N=9 EP=7 IP=8 FDC=26
M0 8 4 3 3 nmos_io_a L=2.8e-07 W=7.4e-05 AD=7.12574e-12 AS=2.21449e-13 PD=3.91524e-06 PS=1.95762e-06 w_cont=2.66e-05 nfing=1 $X=620 $Y=103920 $D=0
X1 1 7 8 9 4 5 3 Usub_7V_ESD $T=0 0 0 0 $X=0 $Y=-3160
.ENDS
***************************************
.SUBCKT ICV_130 1 3 4 5 7 8 9
** N=9 EP=7 IP=8 FDC=26
M0 8 4 3 3 nmos_io_a L=2.8e-07 W=7.4e-05 AD=7.12574e-12 AS=2.21449e-13 PD=3.91524e-06 PS=1.95762e-06 w_cont=2.66e-05 nfing=1 $X=620 $Y=103920 $D=0
X1 1 7 8 9 4 5 3 Usub_7V_ESD $T=0 0 0 0 $X=0 $Y=-3160
.ENDS
***************************************
.SUBCKT ICV_131 1 3 4 5 7 8 9
** N=9 EP=7 IP=8 FDC=26
M0 8 4 3 3 nmos_io_a L=2.8e-07 W=7.4e-05 AD=7.12574e-12 AS=2.21449e-13 PD=3.91524e-06 PS=1.95762e-06 w_cont=2.66e-05 nfing=1 $X=620 $Y=103920 $D=0
X1 1 7 8 9 4 5 3 Usub_7V_ESD $T=0 0 0 0 $X=0 $Y=-3160
.ENDS
***************************************
.SUBCKT ICV_132 1 3 4 5 7 8 9
** N=9 EP=7 IP=8 FDC=26
M0 8 4 3 3 nmos_io_a L=2.8e-07 W=7.4e-05 AD=7.12574e-12 AS=2.21449e-13 PD=3.91524e-06 PS=1.95762e-06 w_cont=2.66e-05 nfing=1 $X=620 $Y=103920 $D=0
X1 1 7 8 9 4 5 3 Usub_7V_ESD $T=0 0 0 0 $X=0 $Y=-3160
.ENDS
***************************************
.SUBCKT nmos_a_CDNS_5887047866546
** N=3 EP=0 IP=0 FDC=0
*.SEEDPROM
.ENDS
***************************************
.SUBCKT ICV_133 1 2 3 4 5 6 7 8 9 10 11 12
** N=17 EP=12 IP=6 FDC=106
*.SEEDPROM
M0 6 5 1 1 nmos_a L=2.4e-07 W=4.8e-07 AD=4.32e-13 AS=2.496e-13 PD=1.08e-06 PS=5.4e-07 w_cont=6e-07 nfing=1 source_num=2 $X=-194480 $Y=272160 $D=1
M1 1 4 1 1 nmos_a L=2e-06 W=5.5e-06 AD=8.30487e-13 AS=1.43e-12 PD=1.59709e-06 PS=1.59709e-06 w_cont=6e-07 nfing=1 source_num=2 $X=-193820 $Y=275380 $D=1
M2 15 7 1 1 nmos_a L=2.4e-07 W=4.8e-07 AD=4.32e-13 AS=2.496e-13 PD=1.08e-06 PS=5.4e-07 w_cont=6e-07 nfing=1 source_num=2 $X=-193720 $Y=272160 $D=1
M3 5 8 15 15 nmos_a L=2.4e-07 W=4.8e-07 AD=4.32e-13 AS=1.92e-13 PD=1.08e-06 PS=5.4e-07 w_cont=6e-07 nfing=1 source_num=2 $X=-192320 $Y=272160 $D=1
M4 1 4 1 1 nmos_a L=2e-06 W=5.5e-06 AD=8.30487e-13 AS=1.43e-12 PD=1.59709e-06 PS=1.59709e-06 w_cont=6e-07 nfing=1 source_num=2 $X=-191300 $Y=275380 $D=1
M5 8 10 1 1 nmos_a L=2.4e-07 W=4.8e-07 AD=4.32e-13 AS=2.496e-13 PD=1.08e-06 PS=5.4e-07 w_cont=6e-07 nfing=1 source_num=2 $X=-190700 $Y=272160 $D=1
M6 10 9 1 1 nmos_a L=4.8e-07 W=4.8e-07 AD=4.32e-13 AS=2.496e-13 PD=1.08e-06 PS=5.4e-07 w_cont=6e-07 nfing=1 source_num=2 $X=-189940 $Y=272160 $D=1
M7 1 4 1 1 nmos_a L=2e-06 W=5.5e-06 AD=8.30487e-13 AS=1.43e-12 PD=1.59709e-06 PS=1.59709e-06 w_cont=6e-07 nfing=1 source_num=2 $X=-188780 $Y=275380 $D=1
M8 10 3 17 17 nmos_a L=4.8e-07 W=4.8e-07 AD=5.832e-13 AS=2.88e-13 PD=1.08e-06 PS=5.4e-07 w_cont=6e-07 nfing=1 source_num=2 $X=-187740 $Y=270140 $D=1
M9 1 4 1 1 nmos_a L=2e-06 W=5.5e-06 AD=8.30487e-13 AS=2.2e-12 PD=1.59709e-06 PS=1.59709e-06 w_cont=6e-07 nfing=1 source_num=2 $X=-186260 $Y=275380 $D=1
M10 12 5 1 1 nmos_a L=2.4e-07 W=1.2e-06 AD=4.68e-13 AS=4.8e-13 PD=9e-07 PS=9e-07 w_cont=6e-07 nfing=1 source_num=2 $X=-185300 $Y=271520 $D=1
M11 12 5 1 1 nmos_a L=2.4e-07 W=1.2e-06 AD=4.68e-13 AS=4.8e-13 PD=9e-07 PS=9e-07 w_cont=6e-07 nfing=1 source_num=2 $X=-184540 $Y=271520 $D=1
M12 1 2 1 1 nmos_a L=2e-06 W=7e-06 AD=8.12983e-13 AS=2.8e-12 PD=1.56343e-06 PS=1.56343e-06 w_cont=6e-07 nfing=1 source_num=2 $X=-182520 $Y=273880 $D=1
M13 1 2 1 1 nmos_a L=2e-06 W=7e-06 AD=8.12983e-13 AS=3.64e-12 PD=1.56343e-06 PS=1.56343e-06 w_cont=6e-07 nfing=1 source_num=2 $X=-180000 $Y=273880 $D=1
M14 1 2 1 1 nmos_a L=2e-06 W=7e-06 AD=8.12983e-13 AS=3.64e-12 PD=1.56343e-06 PS=1.56343e-06 w_cont=6e-07 nfing=1 source_num=2 $X=-177480 $Y=273880 $D=1
M15 1 2 1 1 nmos_a L=2e-06 W=7e-06 AD=8.12983e-13 AS=3.64e-12 PD=1.56343e-06 PS=1.56343e-06 w_cont=6e-07 nfing=1 source_num=2 $X=-174960 $Y=273880 $D=1
M16 1 2 1 1 nmos_a L=2e-06 W=7e-06 AD=8.12983e-13 AS=3.64e-12 PD=1.56343e-06 PS=1.56343e-06 w_cont=6e-07 nfing=1 source_num=2 $X=-172440 $Y=273880 $D=1
M17 1 2 1 1 nmos_a L=2e-06 W=7e-06 AD=8.12983e-13 AS=3.64e-12 PD=1.56343e-06 PS=1.56343e-06 w_cont=6e-07 nfing=1 source_num=2 $X=-169920 $Y=273880 $D=1
M18 1 2 1 1 nmos_a L=2e-06 W=7e-06 AD=8.12983e-13 AS=3.64e-12 PD=1.56343e-06 PS=1.56343e-06 w_cont=6e-07 nfing=1 source_num=2 $X=-167400 $Y=273880 $D=1
M19 1 2 1 1 nmos_a L=2e-06 W=7e-06 AD=8.12983e-13 AS=3.64e-12 PD=1.56343e-06 PS=1.56343e-06 w_cont=6e-07 nfing=1 source_num=2 $X=-164880 $Y=273880 $D=1
M20 1 2 1 1 nmos_a L=2e-06 W=7e-06 AD=8.12983e-13 AS=3.64e-12 PD=1.56343e-06 PS=1.56343e-06 w_cont=6e-07 nfing=1 source_num=2 $X=-162360 $Y=273880 $D=1
M21 1 2 1 1 nmos_a L=2e-06 W=7e-06 AD=8.12983e-13 AS=3.64e-12 PD=1.56343e-06 PS=1.56343e-06 w_cont=6e-07 nfing=1 source_num=2 $X=-159840 $Y=273880 $D=1
M22 1 2 1 1 nmos_a L=2e-06 W=7e-06 AD=8.12983e-13 AS=3.64e-12 PD=1.56343e-06 PS=1.56343e-06 w_cont=6e-07 nfing=1 source_num=2 $X=-157320 $Y=273880 $D=1
M23 1 2 1 1 nmos_a L=2e-06 W=7e-06 AD=8.12983e-13 AS=3.64e-12 PD=1.56343e-06 PS=1.56343e-06 w_cont=6e-07 nfing=1 source_num=2 $X=-154800 $Y=273880 $D=1
M24 1 2 1 1 nmos_a L=2e-06 W=7e-06 AD=8.12983e-13 AS=3.64e-12 PD=1.56343e-06 PS=1.56343e-06 w_cont=6e-07 nfing=1 source_num=2 $X=-152280 $Y=273880 $D=1
M25 1 2 1 1 nmos_a L=2e-06 W=7e-06 AD=8.12983e-13 AS=3.64e-12 PD=1.56343e-06 PS=1.56343e-06 w_cont=6e-07 nfing=1 source_num=2 $X=-149760 $Y=273880 $D=1
M26 1 2 1 1 nmos_a L=2e-06 W=7e-06 AD=8.12983e-13 AS=3.64e-12 PD=1.56343e-06 PS=1.56343e-06 w_cont=6e-07 nfing=1 source_num=2 $X=-147240 $Y=273880 $D=1
M27 1 2 1 1 nmos_a L=2e-06 W=7e-06 AD=8.12983e-13 AS=3.64e-12 PD=1.56343e-06 PS=1.56343e-06 w_cont=6e-07 nfing=1 source_num=2 $X=-144720 $Y=273880 $D=1
M28 1 2 1 1 nmos_a L=2e-06 W=7e-06 AD=8.12983e-13 AS=3.64e-12 PD=1.56343e-06 PS=1.56343e-06 w_cont=6e-07 nfing=1 source_num=2 $X=-142200 $Y=273880 $D=1
M29 1 2 1 1 nmos_a L=2e-06 W=7e-06 AD=8.12983e-13 AS=3.64e-12 PD=1.56343e-06 PS=1.56343e-06 w_cont=6e-07 nfing=1 source_num=2 $X=-139680 $Y=273880 $D=1
M30 1 2 1 1 nmos_a L=2e-06 W=7e-06 AD=8.12983e-13 AS=3.64e-12 PD=1.56343e-06 PS=1.56343e-06 w_cont=6e-07 nfing=1 source_num=2 $X=-137160 $Y=273880 $D=1
M31 1 2 1 1 nmos_a L=2e-06 W=7e-06 AD=8.12983e-13 AS=3.64e-12 PD=1.56343e-06 PS=1.56343e-06 w_cont=6e-07 nfing=1 source_num=2 $X=-134640 $Y=273880 $D=1
M32 1 2 1 1 nmos_a L=2e-06 W=7e-06 AD=8.12983e-13 AS=3.64e-12 PD=1.56343e-06 PS=1.56343e-06 w_cont=6e-07 nfing=1 source_num=2 $X=-132120 $Y=273880 $D=1
M33 1 2 1 1 nmos_a L=2e-06 W=7e-06 AD=8.12983e-13 AS=3.64e-12 PD=1.56343e-06 PS=1.56343e-06 w_cont=6e-07 nfing=1 source_num=2 $X=-129600 $Y=273880 $D=1
M34 1 2 1 1 nmos_a L=2e-06 W=7e-06 AD=8.12983e-13 AS=3.64e-12 PD=1.56343e-06 PS=1.56343e-06 w_cont=6e-07 nfing=1 source_num=2 $X=-127080 $Y=273880 $D=1
M35 1 2 1 1 nmos_a L=2e-06 W=7e-06 AD=8.12983e-13 AS=3.64e-12 PD=1.56343e-06 PS=1.56343e-06 w_cont=6e-07 nfing=1 source_num=2 $X=-124560 $Y=273880 $D=1
M36 1 2 1 1 nmos_a L=2e-06 W=7e-06 AD=8.12983e-13 AS=3.64e-12 PD=1.56343e-06 PS=1.56343e-06 w_cont=6e-07 nfing=1 source_num=2 $X=-122040 $Y=273880 $D=1
M37 1 2 1 1 nmos_a L=2e-06 W=7e-06 AD=8.12983e-13 AS=3.64e-12 PD=1.56343e-06 PS=1.56343e-06 w_cont=6e-07 nfing=1 source_num=2 $X=-119520 $Y=273880 $D=1
M38 1 2 1 1 nmos_a L=2e-06 W=7e-06 AD=8.12983e-13 AS=3.64e-12 PD=1.56343e-06 PS=1.56343e-06 w_cont=6e-07 nfing=1 source_num=2 $X=-117000 $Y=273880 $D=1
M39 1 2 1 1 nmos_a L=2e-06 W=7e-06 AD=8.12983e-13 AS=3.64e-12 PD=1.56343e-06 PS=1.56343e-06 w_cont=6e-07 nfing=1 source_num=2 $X=-114480 $Y=273880 $D=1
M40 1 2 1 1 nmos_a L=2e-06 W=7e-06 AD=8.12983e-13 AS=3.64e-12 PD=1.56343e-06 PS=1.56343e-06 w_cont=6e-07 nfing=1 source_num=2 $X=-111960 $Y=273880 $D=1
M41 1 2 1 1 nmos_a L=2e-06 W=7e-06 AD=8.12983e-13 AS=3.64e-12 PD=1.56343e-06 PS=1.56343e-06 w_cont=6e-07 nfing=1 source_num=2 $X=-109440 $Y=273880 $D=1
M42 1 2 1 1 nmos_a L=2e-06 W=7e-06 AD=8.12983e-13 AS=3.64e-12 PD=1.56343e-06 PS=1.56343e-06 w_cont=6e-07 nfing=1 source_num=2 $X=-106920 $Y=273880 $D=1
M43 1 2 1 1 nmos_a L=2e-06 W=7e-06 AD=8.12983e-13 AS=3.64e-12 PD=1.56343e-06 PS=1.56343e-06 w_cont=6e-07 nfing=1 source_num=2 $X=-104400 $Y=273880 $D=1
M44 1 2 1 1 nmos_a L=2e-06 W=7e-06 AD=8.12983e-13 AS=3.64e-12 PD=1.56343e-06 PS=1.56343e-06 w_cont=6e-07 nfing=1 source_num=2 $X=-101880 $Y=273880 $D=1
M45 1 2 1 1 nmos_a L=2e-06 W=7e-06 AD=8.12983e-13 AS=3.64e-12 PD=1.56343e-06 PS=1.56343e-06 w_cont=6e-07 nfing=1 source_num=2 $X=-99360 $Y=273880 $D=1
M46 1 2 1 1 nmos_a L=2e-06 W=7e-06 AD=8.12983e-13 AS=3.64e-12 PD=1.56343e-06 PS=1.56343e-06 w_cont=6e-07 nfing=1 source_num=2 $X=-96840 $Y=273880 $D=1
M47 1 2 1 1 nmos_a L=2e-06 W=7e-06 AD=8.12983e-13 AS=3.64e-12 PD=1.56343e-06 PS=1.56343e-06 w_cont=6e-07 nfing=1 source_num=2 $X=-94320 $Y=273880 $D=1
M48 1 2 1 1 nmos_a L=2e-06 W=7e-06 AD=8.12983e-13 AS=3.64e-12 PD=1.56343e-06 PS=1.56343e-06 w_cont=6e-07 nfing=1 source_num=2 $X=-91800 $Y=273880 $D=1
M49 1 2 1 1 nmos_a L=2e-06 W=7e-06 AD=8.12983e-13 AS=3.64e-12 PD=1.56343e-06 PS=1.56343e-06 w_cont=6e-07 nfing=1 source_num=2 $X=-89280 $Y=273880 $D=1
M50 1 2 1 1 nmos_a L=2e-06 W=7e-06 AD=8.12983e-13 AS=3.64e-12 PD=1.56343e-06 PS=1.56343e-06 w_cont=6e-07 nfing=1 source_num=2 $X=-86760 $Y=273880 $D=1
M51 1 2 1 1 nmos_a L=2e-06 W=7e-06 AD=8.12983e-13 AS=3.64e-12 PD=1.56343e-06 PS=1.56343e-06 w_cont=6e-07 nfing=1 source_num=2 $X=-84240 $Y=273880 $D=1
M52 1 2 1 1 nmos_a L=2e-06 W=7e-06 AD=8.12983e-13 AS=3.64e-12 PD=1.56343e-06 PS=1.56343e-06 w_cont=6e-07 nfing=1 source_num=2 $X=-81720 $Y=273880 $D=1
M53 1 2 1 1 nmos_a L=2e-06 W=7e-06 AD=8.12983e-13 AS=2.8e-12 PD=1.56343e-06 PS=1.56343e-06 w_cont=6e-07 nfing=1 source_num=2 $X=-79200 $Y=273880 $D=1
M54 11 4 9 9 nmos_a L=3e-07 W=1.2e-06 AD=7.2e-13 AS=4.8e-13 PD=1.8e-06 PS=9e-07 w_cont=6e-07 nfing=1 source_num=2 $X=-188260 $Y=272200 $D=1
M55 17 4 1 1 nmos_a L=3e-07 W=1.2e-06 AD=7.2e-13 AS=4.8e-13 PD=1.8e-06 PS=9e-07 w_cont=6e-07 nfing=1 source_num=2 $X=-186800 $Y=272200 $D=1
M56 16 11 2 2 pmos_a L=2.4e-07 W=4.8e-07 AD=4.32e-13 AS=1.224e-13 PD=1.08e-06 PS=5.4e-07 w_cont=6e-07 nfing=1 mmm=1 $X=-189940 $Y=269000 $D=5
M57 10 3 16 16 pmos_a L=2.4e-07 W=4.8e-07 AD=4.32e-13 AS=1.584e-13 PD=1.08e-06 PS=5.4e-07 w_cont=6e-07 nfing=1 mmm=1 $X=-189940 $Y=270380 $D=5
M58 10 8 16 16 pmos_a L=2.4e-07 W=4.8e-07 AD=4.32e-13 AS=1.584e-13 PD=1.08e-06 PS=5.4e-07 w_cont=6e-07 nfing=1 mmm=1 $X=-189940 $Y=271140 $D=5
M59 2 1 2 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=-194280 $Y=283540 $D=22
M60 2 1 2 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=-191760 $Y=283540 $D=22
M61 2 1 2 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=-189240 $Y=283540 $D=22
M62 2 1 2 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=-186720 $Y=283540 $D=22
M63 2 1 2 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=-184200 $Y=283540 $D=22
M64 2 1 2 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=-181680 $Y=283540 $D=22
M65 2 1 2 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=-179160 $Y=283540 $D=22
M66 2 1 2 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=-176640 $Y=283540 $D=22
M67 2 1 2 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=-174120 $Y=283540 $D=22
M68 2 1 2 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=-171600 $Y=283540 $D=22
M69 2 1 2 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=-169080 $Y=283540 $D=22
M70 2 1 2 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=-166560 $Y=283540 $D=22
M71 2 1 2 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=-164040 $Y=283540 $D=22
M72 2 1 2 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=-161520 $Y=283540 $D=22
M73 2 1 2 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=-159000 $Y=283540 $D=22
M74 2 1 2 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=-156480 $Y=283540 $D=22
M75 2 1 2 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=-153960 $Y=283540 $D=22
M76 2 1 2 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=-151440 $Y=283540 $D=22
M77 2 1 2 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=-148920 $Y=283540 $D=22
M78 2 1 2 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=-146400 $Y=283540 $D=22
M79 2 1 2 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=-143880 $Y=283540 $D=22
M80 2 1 2 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=-141360 $Y=283540 $D=22
M81 2 1 2 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=-138840 $Y=283540 $D=22
M82 2 1 2 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=-136320 $Y=283540 $D=22
M83 2 1 2 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=-133800 $Y=283540 $D=22
M84 2 1 2 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=-131280 $Y=283540 $D=22
M85 2 1 2 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=-128760 $Y=283540 $D=22
M86 2 1 2 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=-126240 $Y=283540 $D=22
M87 2 1 2 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=-123720 $Y=283540 $D=22
M88 2 1 2 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=-121200 $Y=283540 $D=22
M89 2 1 2 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=-118680 $Y=283540 $D=22
M90 2 1 2 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=-116160 $Y=283540 $D=22
M91 2 1 2 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=-113640 $Y=283540 $D=22
M92 2 1 2 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=-111120 $Y=283540 $D=22
M93 2 1 2 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=-108600 $Y=283540 $D=22
M94 2 1 2 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=-106080 $Y=283540 $D=22
M95 2 1 2 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=-103560 $Y=283540 $D=22
M96 2 1 2 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=-101040 $Y=283540 $D=22
M97 2 1 2 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=-98520 $Y=283540 $D=22
M98 2 1 2 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=-96000 $Y=283540 $D=22
M99 2 1 2 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=-93480 $Y=283540 $D=22
M100 2 1 2 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=-90960 $Y=283540 $D=22
M101 2 1 2 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=-88440 $Y=283540 $D=22
M102 2 1 2 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=-85920 $Y=283540 $D=22
M103 2 1 2 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=-83400 $Y=283540 $D=22
M104 2 1 2 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=-80880 $Y=283540 $D=22
M105 2 1 2 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=1.67141e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=-78360 $Y=283540 $D=22
.ENDS
***************************************
.SUBCKT nmos_a_CDNS_5887047866555
** N=2 EP=0 IP=0 FDC=0
*.SEEDPROM
.ENDS
***************************************
.SUBCKT ICV_134
** N=2 EP=0 IP=4 FDC=0
*.SEEDPROM
.ENDS
***************************************
.SUBCKT ICV_135 1 2
** N=2 EP=2 IP=4 FDC=3
*.SEEDPROM
M0 1 2 1 1 nmos_a L=2e-06 W=9.26e-05 AD=7.90041e-13 AS=2.4076e-11 PD=1.51931e-06 PS=1.51931e-06 w_cont=5.1e-06 nfing=1 source_num=2 $X=3140 $Y=200 $D=1
M1 1 2 1 1 nmos_a L=2e-06 W=9.26e-05 AD=7.90041e-13 AS=2.4076e-11 PD=1.51931e-06 PS=1.51931e-06 w_cont=5.1e-06 nfing=1 source_num=2 $X=5660 $Y=200 $D=1
M2 1 2 1 1 nmos_a L=2e-06 W=9.26e-05 AD=7.90041e-13 AS=2.4076e-11 PD=1.51931e-06 PS=1.51931e-06 w_cont=5.1e-06 nfing=1 source_num=2 $X=8180 $Y=200 $D=1
.ENDS
***************************************
.SUBCKT pmos_a_CDNS_5887047866552 1 2 3
** N=3 EP=3 IP=0 FDC=1
M0 2 3 1 1 pmos_a L=2.4e-07 W=9.6e-06 AD=2.568e-12 AS=1.608e-13 PD=6.42e-06 PS=3.21e-06 w_cont=1.1e-06 nfing=1 mmm=1 $X=620 $Y=200 $D=5
.ENDS
***************************************
.SUBCKT pmos_a_CDNS_5887047866541 1 2
** N=2 EP=2 IP=0 FDC=1
M0 1 2 1 1 pmos_a L=2e-06 W=1e-06 AD=6.4e-13 AS=1.25e-13 PD=1.6e-06 PS=8e-07 w_cont=6e-07 nfing=1 mmm=1 $X=620 $Y=200 $D=5
.ENDS
***************************************
.SUBCKT ICV_136 1 2 4 8 9 10 12
** N=13 EP=7 IP=56 FDC=59
*.SEEDPROM
M0 4 12 4 4 nmos_a L=2e-06 W=9.26e-05 AD=7.90041e-13 AS=2.4076e-11 PD=1.51931e-06 PS=1.51931e-06 w_cont=5.1e-06 nfing=1 source_num=2 $X=-81620 $Y=160080 $D=1
M1 4 12 4 4 nmos_a L=2e-06 W=9.26e-05 AD=7.90041e-13 AS=3.704e-11 PD=1.51931e-06 PS=1.51931e-06 w_cont=5.1e-06 nfing=1 source_num=2 $X=-79100 $Y=160080 $D=1
M2 4 12 4 4 nmos_a L=2e-06 W=9.26e-05 AD=7.90041e-13 AS=3.704e-11 PD=1.51931e-06 PS=1.51931e-06 w_cont=5.1e-06 nfing=1 source_num=2 $X=-192500 $Y=160080 $D=1
M3 4 12 4 4 nmos_a L=2e-06 W=9.26e-05 AD=7.90041e-13 AS=2.4076e-11 PD=1.51931e-06 PS=1.51931e-06 w_cont=5.1e-06 nfing=1 source_num=2 $X=-182420 $Y=160080 $D=1
M4 4 12 4 4 nmos_a L=2e-06 W=9.26e-05 AD=7.90041e-13 AS=2.4076e-11 PD=1.51931e-06 PS=1.51931e-06 w_cont=5.1e-06 nfing=1 source_num=2 $X=-172340 $Y=160080 $D=1
M5 4 12 4 4 nmos_a L=2e-06 W=9.26e-05 AD=7.90041e-13 AS=2.4076e-11 PD=1.51931e-06 PS=1.51931e-06 w_cont=5.1e-06 nfing=1 source_num=2 $X=-162260 $Y=160080 $D=1
M6 4 12 4 4 nmos_a L=2e-06 W=9.26e-05 AD=7.90041e-13 AS=2.4076e-11 PD=1.51931e-06 PS=1.51931e-06 w_cont=5.1e-06 nfing=1 source_num=2 $X=-152180 $Y=160080 $D=1
M7 4 12 4 4 nmos_a L=2e-06 W=9.26e-05 AD=7.90041e-13 AS=2.4076e-11 PD=1.51931e-06 PS=1.51931e-06 w_cont=5.1e-06 nfing=1 source_num=2 $X=-142100 $Y=160080 $D=1
M8 4 12 4 4 nmos_a L=2e-06 W=9.26e-05 AD=7.90041e-13 AS=2.4076e-11 PD=1.51931e-06 PS=1.51931e-06 w_cont=5.1e-06 nfing=1 source_num=2 $X=-132020 $Y=160080 $D=1
M9 4 12 4 4 nmos_a L=2e-06 W=9.26e-05 AD=7.90041e-13 AS=2.4076e-11 PD=1.51931e-06 PS=1.51931e-06 w_cont=5.1e-06 nfing=1 source_num=2 $X=-121940 $Y=160080 $D=1
M10 4 12 4 4 nmos_a L=2e-06 W=9.26e-05 AD=7.90041e-13 AS=2.4076e-11 PD=1.51931e-06 PS=1.51931e-06 w_cont=5.1e-06 nfing=1 source_num=2 $X=-111860 $Y=160080 $D=1
M11 4 12 4 4 nmos_a L=2e-06 W=9.26e-05 AD=7.90041e-13 AS=2.4076e-11 PD=1.51931e-06 PS=1.51931e-06 w_cont=5.1e-06 nfing=1 source_num=2 $X=-101780 $Y=160080 $D=1
M12 4 12 4 4 nmos_a L=2e-06 W=9.26e-05 AD=7.90041e-13 AS=2.4076e-11 PD=1.51931e-06 PS=1.51931e-06 w_cont=5.1e-06 nfing=1 source_num=2 $X=-91700 $Y=160080 $D=1
M13 8 10 2 2 pmos_a L=2.4e-07 W=4.8e-07 AD=4.32e-13 AS=1.224e-13 PD=1.08e-06 PS=5.4e-07 w_cont=6e-07 nfing=1 mmm=1 $X=-189920 $Y=267560 $D=5
M14 9 10 2 2 pmos_a L=2.4e-07 W=4.8e-07 AD=4.32e-13 AS=1.224e-13 PD=1.08e-06 PS=5.4e-07 w_cont=6e-07 nfing=1 mmm=1 $X=-188440 $Y=267560 $D=5
X15 1 4 10 nmos_a_CDNS_5887047866553 $T=-169060 259920 0 270 $X=-169060 $Y=258480
X16 1 4 10 nmos_a_CDNS_5887047866553 $T=-149660 259920 0 270 $X=-149660 $Y=258480
X17 1 4 10 nmos_a_CDNS_5887047866553 $T=-130100 259920 0 270 $X=-130100 $Y=258480
X18 1 4 10 nmos_a_CDNS_5887047866553 $T=-110700 259920 0 270 $X=-110700 $Y=258480
X19 1 4 10 nmos_a_CDNS_5887047866553 $T=-91300 259920 0 270 $X=-91300 $Y=258480
X21 4 12 ICV_135 $T=-193120 159880 0 0 $X=-193120 $Y=159880
X22 4 12 ICV_135 $T=-183040 159880 0 0 $X=-183040 $Y=159880
X23 4 12 ICV_135 $T=-172960 159880 0 0 $X=-172960 $Y=159880
X24 4 12 ICV_135 $T=-162880 159880 0 0 $X=-162880 $Y=159880
X25 4 12 ICV_135 $T=-152800 159880 0 0 $X=-152800 $Y=159880
X26 4 12 ICV_135 $T=-142720 159880 0 0 $X=-142720 $Y=159880
X27 4 12 ICV_135 $T=-132640 159880 0 0 $X=-132640 $Y=159880
X28 4 12 ICV_135 $T=-122560 159880 0 0 $X=-122560 $Y=159880
X29 4 12 ICV_135 $T=-112480 159880 0 0 $X=-112480 $Y=159880
X30 4 12 ICV_135 $T=-102400 159880 0 0 $X=-102400 $Y=159880
X31 4 12 ICV_135 $T=-92320 159880 0 0 $X=-92320 $Y=159880
X32 2 4 10 pmos_a_CDNS_5887047866552 $T=-169740 258480 0 90 $X=-180840 $Y=258480
X33 2 4 10 pmos_a_CDNS_5887047866552 $T=-150160 258480 0 90 $X=-161260 $Y=258480
X34 2 4 10 pmos_a_CDNS_5887047866552 $T=-130760 258480 0 90 $X=-141860 $Y=258480
X35 2 4 10 pmos_a_CDNS_5887047866552 $T=-111200 258480 0 90 $X=-122300 $Y=258480
X36 2 4 10 pmos_a_CDNS_5887047866552 $T=-91800 258480 0 90 $X=-102900 $Y=258480
X37 2 9 pmos_a_CDNS_5887047866541 $T=-184940 264940 1 180 $X=-188140 $Y=264940
.ENDS
***************************************
.SUBCKT ICV_137
** N=2 EP=0 IP=4 FDC=0
*.SEEDPROM
.ENDS
***************************************
.SUBCKT ICV_138 1 2
** N=2 EP=2 IP=4 FDC=3
*.SEEDPROM
M0 1 2 1 1 nmos_a L=2e-06 W=9.26e-05 AD=7.90041e-13 AS=2.4076e-11 PD=1.51931e-06 PS=1.51931e-06 w_cont=5.1e-06 nfing=1 source_num=2 $X=-6940 $Y=200 $D=1
M1 1 2 1 1 nmos_a L=2e-06 W=9.26e-05 AD=7.90041e-13 AS=2.4076e-11 PD=1.51931e-06 PS=1.51931e-06 w_cont=5.1e-06 nfing=1 source_num=2 $X=-4420 $Y=200 $D=1
M2 1 2 1 1 nmos_a L=2e-06 W=9.26e-05 AD=7.90041e-13 AS=2.4076e-11 PD=1.51931e-06 PS=1.51931e-06 w_cont=5.1e-06 nfing=1 source_num=2 $X=-1900 $Y=200 $D=1
.ENDS
***************************************
.SUBCKT ICV_139 2 3
** N=3 EP=2 IP=24 FDC=46
M0 2 3 2 2 nmos_a L=2e-06 W=9.26e-05 AD=1.21545e-12 AS=2.4076e-11 PD=3.03862e-06 PS=1.51931e-06 w_cont=5.1e-06 nfing=1 source_num=2 $X=-79100 $Y=61480 $D=1
M1 2 3 2 2 nmos_a L=2e-06 W=9.26e-05 AD=7.90041e-13 AS=2.4076e-11 PD=1.51931e-06 PS=1.51931e-06 w_cont=5.1e-06 nfing=1 source_num=2 $X=-81620 $Y=61480 $D=1
M2 2 3 2 2 nmos_a L=2e-06 W=9.26e-05 AD=1.21545e-12 AS=2.4076e-11 PD=3.03862e-06 PS=1.51931e-06 w_cont=5.1e-06 nfing=1 source_num=2 $X=-192500 $Y=61480 $D=1
M3 2 3 2 2 nmos_a L=2e-06 W=9.26e-05 AD=7.90041e-13 AS=2.4076e-11 PD=1.51931e-06 PS=1.51931e-06 w_cont=5.1e-06 nfing=1 source_num=2 $X=-182420 $Y=61480 $D=1
M4 2 3 2 2 nmos_a L=2e-06 W=9.26e-05 AD=7.90041e-13 AS=2.4076e-11 PD=1.51931e-06 PS=1.51931e-06 w_cont=5.1e-06 nfing=1 source_num=2 $X=-172340 $Y=61480 $D=1
M5 2 3 2 2 nmos_a L=2e-06 W=9.26e-05 AD=7.90041e-13 AS=2.4076e-11 PD=1.51931e-06 PS=1.51931e-06 w_cont=5.1e-06 nfing=1 source_num=2 $X=-162260 $Y=61480 $D=1
M6 2 3 2 2 nmos_a L=2e-06 W=9.26e-05 AD=7.90041e-13 AS=2.4076e-11 PD=1.51931e-06 PS=1.51931e-06 w_cont=5.1e-06 nfing=1 source_num=2 $X=-152180 $Y=61480 $D=1
M7 2 3 2 2 nmos_a L=2e-06 W=9.26e-05 AD=7.90041e-13 AS=2.4076e-11 PD=1.51931e-06 PS=1.51931e-06 w_cont=5.1e-06 nfing=1 source_num=2 $X=-142100 $Y=61480 $D=1
M8 2 3 2 2 nmos_a L=2e-06 W=9.26e-05 AD=7.90041e-13 AS=2.4076e-11 PD=1.51931e-06 PS=1.51931e-06 w_cont=5.1e-06 nfing=1 source_num=2 $X=-132020 $Y=61480 $D=1
M9 2 3 2 2 nmos_a L=2e-06 W=9.26e-05 AD=7.90041e-13 AS=2.4076e-11 PD=1.51931e-06 PS=1.51931e-06 w_cont=5.1e-06 nfing=1 source_num=2 $X=-121940 $Y=61480 $D=1
M10 2 3 2 2 nmos_a L=2e-06 W=9.26e-05 AD=7.90041e-13 AS=2.4076e-11 PD=1.51931e-06 PS=1.51931e-06 w_cont=5.1e-06 nfing=1 source_num=2 $X=-111860 $Y=61480 $D=1
M11 2 3 2 2 nmos_a L=2e-06 W=9.26e-05 AD=7.90041e-13 AS=2.4076e-11 PD=1.51931e-06 PS=1.51931e-06 w_cont=5.1e-06 nfing=1 source_num=2 $X=-101780 $Y=61480 $D=1
M12 2 3 2 2 nmos_a L=2e-06 W=9.26e-05 AD=7.90041e-13 AS=2.4076e-11 PD=1.51931e-06 PS=1.51931e-06 w_cont=5.1e-06 nfing=1 source_num=2 $X=-91700 $Y=61480 $D=1
X14 2 3 ICV_138 $T=-189880 61280 1 180 $X=-193080 $Y=61280
X15 2 3 ICV_138 $T=-179800 61280 1 180 $X=-183000 $Y=61280
X16 2 3 ICV_138 $T=-169720 61280 1 180 $X=-172920 $Y=61280
X17 2 3 ICV_138 $T=-159640 61280 1 180 $X=-162840 $Y=61280
X18 2 3 ICV_138 $T=-149560 61280 1 180 $X=-152760 $Y=61280
X19 2 3 ICV_138 $T=-139480 61280 1 180 $X=-142680 $Y=61280
X20 2 3 ICV_138 $T=-129400 61280 1 180 $X=-132600 $Y=61280
X21 2 3 ICV_138 $T=-119320 61280 1 180 $X=-122520 $Y=61280
X22 2 3 ICV_138 $T=-109240 61280 1 180 $X=-112440 $Y=61280
X23 2 3 ICV_138 $T=-99160 61280 1 180 $X=-102360 $Y=61280
X24 2 3 ICV_138 $T=-89080 61280 1 180 $X=-92280 $Y=61280
.ENDS
***************************************
.SUBCKT nmos_a_CDNS_5887047866556
** N=2 EP=0 IP=0 FDC=0
*.SEEDPROM
.ENDS
***************************************
.SUBCKT ICV_140
** N=2 EP=0 IP=4 FDC=0
*.SEEDPROM
.ENDS
***************************************
.SUBCKT nmos_a_CDNS_5887047866550
** N=2 EP=0 IP=0 FDC=0
*.SEEDPROM
.ENDS
***************************************
.SUBCKT ICV_141
** N=2 EP=0 IP=4 FDC=0
*.SEEDPROM
.ENDS
***************************************
.SUBCKT ICV_142 1 2
** N=2 EP=2 IP=4 FDC=3
*.SEEDPROM
M0 1 2 1 1 nmos_a L=2e-06 W=7e-05 AD=7.8731e-13 AS=1.82e-11 PD=1.51406e-06 PS=1.51406e-06 w_cont=3.6e-06 nfing=1 source_num=2 $X=-6940 $Y=200 $D=1
M1 1 2 1 1 nmos_a L=2e-06 W=7e-05 AD=7.8731e-13 AS=1.82e-11 PD=1.51406e-06 PS=1.51406e-06 w_cont=3.6e-06 nfing=1 source_num=2 $X=-4420 $Y=200 $D=1
M2 1 2 1 1 nmos_a L=2e-06 W=7e-05 AD=7.8731e-13 AS=1.82e-11 PD=1.51406e-06 PS=1.51406e-06 w_cont=3.6e-06 nfing=1 source_num=2 $X=-1900 $Y=200 $D=1
.ENDS
***************************************
.SUBCKT ICV_143 1 2
** N=2 EP=2 IP=4 FDC=3
*.SEEDPROM
M0 1 2 1 1 nmos_a L=2e-06 W=1.5e-05 AD=8.03712e-13 AS=3.9e-12 PD=1.5456e-06 PS=1.5456e-06 w_cont=1.1e-06 nfing=1 source_num=2 $X=-6940 $Y=200 $D=1
M1 1 2 1 1 nmos_a L=2e-06 W=1.5e-05 AD=8.03712e-13 AS=3.9e-12 PD=1.5456e-06 PS=1.5456e-06 w_cont=1.1e-06 nfing=1 source_num=2 $X=-4420 $Y=200 $D=1
M2 1 2 1 1 nmos_a L=2e-06 W=1.5e-05 AD=8.03712e-13 AS=3.9e-12 PD=1.5456e-06 PS=1.5456e-06 w_cont=1.1e-06 nfing=1 source_num=2 $X=-1900 $Y=200 $D=1
.ENDS
***************************************
.SUBCKT nmos_a_CDNS_5887047866558 1 2 3
** N=3 EP=3 IP=0 FDC=1
M0 2 3 1 1 nmos_a L=2.8e-07 W=2.4e-06 AD=1.4e-12 AS=9.6e-13 PD=3.5e-06 PS=1.75e-06 w_cont=1.1e-06 nfing=1 source_num=2 $X=620 $Y=200 $D=1
.ENDS
***************************************
.SUBCKT pmos_a_CDNS_5887047866557 1 2 3
** N=3 EP=3 IP=0 FDC=1
M0 2 3 1 1 pmos_a L=2.4e-07 W=4.8e-06 AD=2.16e-12 AS=1.44e-13 PD=5.4e-06 PS=2.7e-06 w_cont=6e-07 nfing=1 mmm=1 $X=620 $Y=200 $D=5
.ENDS
***************************************
.SUBCKT ICV_144 2 3 4 6 7 8 9 10 11 12
** N=12 EP=10 IP=72 FDC=100
M0 12 8 12 12 nmos_a L=2e-06 W=7e-05 AD=1.21125e-12 AS=1.82e-11 PD=3.02811e-06 PS=1.51406e-06 w_cont=3.6e-06 nfing=1 source_num=2 $X=-79100 $Y=-15340 $D=1
M1 12 8 12 12 nmos_a L=2e-06 W=7e-05 AD=7.8731e-13 AS=1.82e-11 PD=1.51406e-06 PS=1.51406e-06 w_cont=3.6e-06 nfing=1 source_num=2 $X=-81620 $Y=-15340 $D=1
M2 11 6 11 11 nmos_a L=2e-06 W=1.5e-05 AD=1.23648e-12 AS=3.9e-12 PD=3.0912e-06 PS=1.5456e-06 w_cont=1.1e-06 nfing=1 source_num=2 $X=-79100 $Y=-34660 $D=1
M3 11 6 11 11 nmos_a L=2e-06 W=1.5e-05 AD=8.03712e-13 AS=3.9e-12 PD=1.5456e-06 PS=1.5456e-06 w_cont=1.1e-06 nfing=1 source_num=2 $X=-81620 $Y=-34660 $D=1
M4 12 8 12 12 nmos_a L=2e-06 W=7e-05 AD=1.21125e-12 AS=1.82e-11 PD=3.02811e-06 PS=1.51406e-06 w_cont=3.6e-06 nfing=1 source_num=2 $X=-192500 $Y=-15340 $D=1
M5 12 8 12 12 nmos_a L=2e-06 W=7e-05 AD=7.8731e-13 AS=1.82e-11 PD=1.51406e-06 PS=1.51406e-06 w_cont=3.6e-06 nfing=1 source_num=2 $X=-182420 $Y=-15340 $D=1
M6 12 8 12 12 nmos_a L=2e-06 W=7e-05 AD=7.8731e-13 AS=1.82e-11 PD=1.51406e-06 PS=1.51406e-06 w_cont=3.6e-06 nfing=1 source_num=2 $X=-172340 $Y=-15340 $D=1
M7 12 8 12 12 nmos_a L=2e-06 W=7e-05 AD=7.8731e-13 AS=1.82e-11 PD=1.51406e-06 PS=1.51406e-06 w_cont=3.6e-06 nfing=1 source_num=2 $X=-162260 $Y=-15340 $D=1
M8 12 8 12 12 nmos_a L=2e-06 W=7e-05 AD=7.8731e-13 AS=1.82e-11 PD=1.51406e-06 PS=1.51406e-06 w_cont=3.6e-06 nfing=1 source_num=2 $X=-152180 $Y=-15340 $D=1
M9 12 8 12 12 nmos_a L=2e-06 W=7e-05 AD=7.8731e-13 AS=1.82e-11 PD=1.51406e-06 PS=1.51406e-06 w_cont=3.6e-06 nfing=1 source_num=2 $X=-142100 $Y=-15340 $D=1
M10 12 8 12 12 nmos_a L=2e-06 W=7e-05 AD=7.8731e-13 AS=1.82e-11 PD=1.51406e-06 PS=1.51406e-06 w_cont=3.6e-06 nfing=1 source_num=2 $X=-132020 $Y=-15340 $D=1
M11 12 8 12 12 nmos_a L=2e-06 W=7e-05 AD=7.8731e-13 AS=1.82e-11 PD=1.51406e-06 PS=1.51406e-06 w_cont=3.6e-06 nfing=1 source_num=2 $X=-121940 $Y=-15340 $D=1
M12 12 8 12 12 nmos_a L=2e-06 W=7e-05 AD=7.8731e-13 AS=1.82e-11 PD=1.51406e-06 PS=1.51406e-06 w_cont=3.6e-06 nfing=1 source_num=2 $X=-111860 $Y=-15340 $D=1
M13 12 8 12 12 nmos_a L=2e-06 W=7e-05 AD=7.8731e-13 AS=1.82e-11 PD=1.51406e-06 PS=1.51406e-06 w_cont=3.6e-06 nfing=1 source_num=2 $X=-101780 $Y=-15340 $D=1
M14 12 8 12 12 nmos_a L=2e-06 W=7e-05 AD=7.8731e-13 AS=1.82e-11 PD=1.51406e-06 PS=1.51406e-06 w_cont=3.6e-06 nfing=1 source_num=2 $X=-91700 $Y=-15340 $D=1
M15 11 6 11 11 nmos_a L=2e-06 W=1.5e-05 AD=1.23648e-12 AS=3.9e-12 PD=3.0912e-06 PS=1.5456e-06 w_cont=1.1e-06 nfing=1 source_num=2 $X=-192500 $Y=-34660 $D=1
M16 11 6 11 11 nmos_a L=2e-06 W=1.5e-05 AD=8.03712e-13 AS=3.9e-12 PD=1.5456e-06 PS=1.5456e-06 w_cont=1.1e-06 nfing=1 source_num=2 $X=-182420 $Y=-34660 $D=1
M17 11 6 11 11 nmos_a L=2e-06 W=1.5e-05 AD=8.03712e-13 AS=3.9e-12 PD=1.5456e-06 PS=1.5456e-06 w_cont=1.1e-06 nfing=1 source_num=2 $X=-172340 $Y=-34660 $D=1
M18 11 6 11 11 nmos_a L=2e-06 W=1.5e-05 AD=8.03712e-13 AS=3.9e-12 PD=1.5456e-06 PS=1.5456e-06 w_cont=1.1e-06 nfing=1 source_num=2 $X=-162260 $Y=-34660 $D=1
M19 11 6 11 11 nmos_a L=2e-06 W=1.5e-05 AD=8.03712e-13 AS=3.9e-12 PD=1.5456e-06 PS=1.5456e-06 w_cont=1.1e-06 nfing=1 source_num=2 $X=-152180 $Y=-34660 $D=1
M20 11 6 11 11 nmos_a L=2e-06 W=1.5e-05 AD=8.03712e-13 AS=3.9e-12 PD=1.5456e-06 PS=1.5456e-06 w_cont=1.1e-06 nfing=1 source_num=2 $X=-142100 $Y=-34660 $D=1
M21 11 6 11 11 nmos_a L=2e-06 W=1.5e-05 AD=8.03712e-13 AS=3.9e-12 PD=1.5456e-06 PS=1.5456e-06 w_cont=1.1e-06 nfing=1 source_num=2 $X=-132020 $Y=-34660 $D=1
M22 11 6 11 11 nmos_a L=2e-06 W=1.5e-05 AD=8.03712e-13 AS=3.9e-12 PD=1.5456e-06 PS=1.5456e-06 w_cont=1.1e-06 nfing=1 source_num=2 $X=-121940 $Y=-34660 $D=1
M23 11 6 11 11 nmos_a L=2e-06 W=1.5e-05 AD=8.03712e-13 AS=3.9e-12 PD=1.5456e-06 PS=1.5456e-06 w_cont=1.1e-06 nfing=1 source_num=2 $X=-111860 $Y=-34660 $D=1
M24 11 6 11 11 nmos_a L=2e-06 W=1.5e-05 AD=8.03712e-13 AS=3.9e-12 PD=1.5456e-06 PS=1.5456e-06 w_cont=1.1e-06 nfing=1 source_num=2 $X=-101780 $Y=-34660 $D=1
M25 11 6 11 11 nmos_a L=2e-06 W=1.5e-05 AD=8.03712e-13 AS=3.9e-12 PD=1.5456e-06 PS=1.5456e-06 w_cont=1.1e-06 nfing=1 source_num=2 $X=-91700 $Y=-34660 $D=1
X26 4 12 7 nmos_a_CDNS_5887047866553 $T=-185200 58960 0 90 $X=-192500 $Y=58960
X27 3 11 8 nmos_a_CDNS_5887047866553 $T=-180400 -17860 1 90 $X=-180400 $Y=-17860
X28 4 12 7 nmos_a_CDNS_5887047866553 $T=-165800 58960 0 90 $X=-173100 $Y=58960
X29 4 11 8 pmos_a_CDNS_5887047866552 $T=-180900 -16380 1 270 $X=-192000 $Y=-17820
X30 2 12 7 pmos_a_CDNS_5887047866552 $T=-184700 60440 0 270 $X=-184700 $Y=59000
X31 2 12 7 pmos_a_CDNS_5887047866552 $T=-165300 60440 0 270 $X=-165300 $Y=59000
X34 12 8 ICV_142 $T=-189880 -15540 1 180 $X=-193080 $Y=-15540
X35 12 8 ICV_142 $T=-179800 -15540 1 180 $X=-183000 $Y=-15540
X36 12 8 ICV_142 $T=-169720 -15540 1 180 $X=-172920 $Y=-15540
X37 12 8 ICV_142 $T=-159640 -15540 1 180 $X=-162840 $Y=-15540
X38 12 8 ICV_142 $T=-149560 -15540 1 180 $X=-152760 $Y=-15540
X39 12 8 ICV_142 $T=-139480 -15540 1 180 $X=-142680 $Y=-15540
X40 12 8 ICV_142 $T=-129400 -15540 1 180 $X=-132600 $Y=-15540
X41 12 8 ICV_142 $T=-119320 -15540 1 180 $X=-122520 $Y=-15540
X42 12 8 ICV_142 $T=-109240 -15540 1 180 $X=-112440 $Y=-15540
X43 12 8 ICV_142 $T=-99160 -15540 1 180 $X=-102360 $Y=-15540
X44 12 8 ICV_142 $T=-89080 -15540 1 180 $X=-92280 $Y=-15540
X45 11 6 ICV_143 $T=-189880 -34860 1 180 $X=-193080 $Y=-34860
X46 11 6 ICV_143 $T=-179800 -34860 1 180 $X=-183000 $Y=-34860
X47 11 6 ICV_143 $T=-169720 -34860 1 180 $X=-172920 $Y=-34860
X48 11 6 ICV_143 $T=-159640 -34860 1 180 $X=-162840 $Y=-34860
X49 11 6 ICV_143 $T=-149560 -34860 1 180 $X=-152760 $Y=-34860
X50 11 6 ICV_143 $T=-139480 -34860 1 180 $X=-142680 $Y=-34860
X51 11 6 ICV_143 $T=-129400 -34860 1 180 $X=-132600 $Y=-34860
X52 11 6 ICV_143 $T=-119320 -34860 1 180 $X=-122520 $Y=-34860
X53 11 6 ICV_143 $T=-109240 -34860 1 180 $X=-112440 $Y=-34860
X54 11 6 ICV_143 $T=-99160 -34860 1 180 $X=-102360 $Y=-34860
X55 11 6 ICV_143 $T=-89080 -34860 1 180 $X=-92280 $Y=-34860
X56 10 9 6 nmos_a_CDNS_5887047866558 $T=-185040 -37180 1 90 $X=-185040 $Y=-37180
X57 3 9 6 pmos_a_CDNS_5887047866557 $T=-185540 -35700 1 270 $X=-191340 $Y=-37140
.ENDS
***************************************
.SUBCKT nmos_a_CDNS_5887047866551
** N=2 EP=0 IP=0 FDC=0
*.SEEDPROM
.ENDS
***************************************
.SUBCKT ICV_145
** N=2 EP=0 IP=4 FDC=0
*.SEEDPROM
.ENDS
***************************************
.SUBCKT ICV_146 1 2
** N=2 EP=2 IP=4 FDC=3
*.SEEDPROM
M0 1 2 1 1 nmos_a L=2e-06 W=0.0001 AD=7.86989e-13 AS=2.6e-11 PD=1.51344e-06 PS=1.51344e-06 w_cont=5.1e-06 nfing=1 source_num=2 $X=-6940 $Y=200 $D=1
M1 1 2 1 1 nmos_a L=2e-06 W=0.0001 AD=7.86989e-13 AS=2.6e-11 PD=1.51344e-06 PS=1.51344e-06 w_cont=5.1e-06 nfing=1 source_num=2 $X=-4420 $Y=200 $D=1
M2 1 2 1 1 nmos_a L=2e-06 W=0.0001 AD=7.86989e-13 AS=2.6e-11 PD=1.51344e-06 PS=1.51344e-06 w_cont=5.1e-06 nfing=1 source_num=2 $X=-1900 $Y=200 $D=1
.ENDS
***************************************
.SUBCKT ICV_147 4 6
** N=7 EP=2 IP=24 FDC=46
M0 4 6 4 4 nmos_a L=2e-06 W=0.0001 AD=1.21075e-12 AS=2.6e-11 PD=3.02688e-06 PS=1.51344e-06 w_cont=5.1e-06 nfing=1 source_num=2 $X=-79100 $Y=-142980 $D=1
M1 4 6 4 4 nmos_a L=2e-06 W=0.0001 AD=7.86989e-13 AS=2.6e-11 PD=1.51344e-06 PS=1.51344e-06 w_cont=5.1e-06 nfing=1 source_num=2 $X=-81620 $Y=-142980 $D=1
M2 4 6 4 4 nmos_a L=2e-06 W=0.0001 AD=1.21075e-12 AS=2.6e-11 PD=3.02688e-06 PS=1.51344e-06 w_cont=5.1e-06 nfing=1 source_num=2 $X=-192500 $Y=-142980 $D=1
M3 4 6 4 4 nmos_a L=2e-06 W=0.0001 AD=7.86989e-13 AS=2.6e-11 PD=1.51344e-06 PS=1.51344e-06 w_cont=5.1e-06 nfing=1 source_num=2 $X=-182420 $Y=-142980 $D=1
M4 4 6 4 4 nmos_a L=2e-06 W=0.0001 AD=7.86989e-13 AS=2.6e-11 PD=1.51344e-06 PS=1.51344e-06 w_cont=5.1e-06 nfing=1 source_num=2 $X=-172340 $Y=-142980 $D=1
M5 4 6 4 4 nmos_a L=2e-06 W=0.0001 AD=7.86989e-13 AS=2.6e-11 PD=1.51344e-06 PS=1.51344e-06 w_cont=5.1e-06 nfing=1 source_num=2 $X=-162260 $Y=-142980 $D=1
M6 4 6 4 4 nmos_a L=2e-06 W=0.0001 AD=7.86989e-13 AS=2.6e-11 PD=1.51344e-06 PS=1.51344e-06 w_cont=5.1e-06 nfing=1 source_num=2 $X=-152180 $Y=-142980 $D=1
M7 4 6 4 4 nmos_a L=2e-06 W=0.0001 AD=7.86989e-13 AS=2.6e-11 PD=1.51344e-06 PS=1.51344e-06 w_cont=5.1e-06 nfing=1 source_num=2 $X=-142100 $Y=-142980 $D=1
M8 4 6 4 4 nmos_a L=2e-06 W=0.0001 AD=7.86989e-13 AS=2.6e-11 PD=1.51344e-06 PS=1.51344e-06 w_cont=5.1e-06 nfing=1 source_num=2 $X=-132020 $Y=-142980 $D=1
M9 4 6 4 4 nmos_a L=2e-06 W=0.0001 AD=7.86989e-13 AS=2.6e-11 PD=1.51344e-06 PS=1.51344e-06 w_cont=5.1e-06 nfing=1 source_num=2 $X=-121940 $Y=-142980 $D=1
M10 4 6 4 4 nmos_a L=2e-06 W=0.0001 AD=7.86989e-13 AS=2.6e-11 PD=1.51344e-06 PS=1.51344e-06 w_cont=5.1e-06 nfing=1 source_num=2 $X=-111860 $Y=-142980 $D=1
M11 4 6 4 4 nmos_a L=2e-06 W=0.0001 AD=7.86989e-13 AS=2.6e-11 PD=1.51344e-06 PS=1.51344e-06 w_cont=5.1e-06 nfing=1 source_num=2 $X=-101780 $Y=-142980 $D=1
M12 4 6 4 4 nmos_a L=2e-06 W=0.0001 AD=7.86989e-13 AS=2.6e-11 PD=1.51344e-06 PS=1.51344e-06 w_cont=5.1e-06 nfing=1 source_num=2 $X=-91700 $Y=-142980 $D=1
X14 4 6 ICV_146 $T=-189880 -143180 1 180 $X=-193080 $Y=-143180
X15 4 6 ICV_146 $T=-179800 -143180 1 180 $X=-183000 $Y=-143180
X16 4 6 ICV_146 $T=-169720 -143180 1 180 $X=-172920 $Y=-143180
X17 4 6 ICV_146 $T=-159640 -143180 1 180 $X=-162840 $Y=-143180
X18 4 6 ICV_146 $T=-149560 -143180 1 180 $X=-152760 $Y=-143180
X19 4 6 ICV_146 $T=-139480 -143180 1 180 $X=-142680 $Y=-143180
X20 4 6 ICV_146 $T=-129400 -143180 1 180 $X=-132600 $Y=-143180
X21 4 6 ICV_146 $T=-119320 -143180 1 180 $X=-122520 $Y=-143180
X22 4 6 ICV_146 $T=-109240 -143180 1 180 $X=-112440 $Y=-143180
X23 4 6 ICV_146 $T=-99160 -143180 1 180 $X=-102360 $Y=-143180
X24 4 6 ICV_146 $T=-89080 -143180 1 180 $X=-92280 $Y=-143180
.ENDS
***************************************
.SUBCKT nmos_a_CDNS_5887047866547 1 2 3
** N=3 EP=3 IP=0 FDC=1
M0 2 3 1 1 nmos_a L=2.4e-07 W=7.2e-06 AD=1.648e-12 AS=2.88e-12 PD=4.12e-06 PS=2.06e-06 w_cont=3.1e-06 nfing=1 source_num=2 $X=620 $Y=200 $D=1
.ENDS
***************************************
.SUBCKT ICV_148 2 3 4 5
** N=21 EP=4 IP=84 FDC=28
*.SEEDPROM
M0 7 7 8 8 nmos_a L=2.4e-07 W=1.2e-06 AD=7.2e-13 AS=4.8e-13 PD=1.8e-06 PS=9e-07 w_cont=6e-07 nfing=1 source_num=2 $X=-188540 $Y=-144820 $D=1
M1 9 9 4 4 nmos_a L=2.4e-07 W=1.2e-06 AD=7.2e-13 AS=4.8e-13 PD=1.8e-06 PS=9e-07 w_cont=6e-07 nfing=1 source_num=2 $X=-183140 $Y=-144820 $D=1
M2 10 10 11 11 nmos_a L=2.4e-07 W=1.2e-06 AD=7.2e-13 AS=4.8e-13 PD=1.8e-06 PS=9e-07 w_cont=6e-07 nfing=1 source_num=2 $X=-163340 $Y=-144820 $D=1
M3 12 12 4 4 nmos_a L=2.4e-07 W=1.2e-06 AD=7.2e-13 AS=4.8e-13 PD=1.8e-06 PS=9e-07 w_cont=6e-07 nfing=1 source_num=2 $X=-157940 $Y=-144820 $D=1
M4 13 13 14 14 nmos_a L=2.4e-07 W=1.2e-06 AD=7.2e-13 AS=4.8e-13 PD=1.8e-06 PS=9e-07 w_cont=6e-07 nfing=1 source_num=2 $X=-138140 $Y=-144820 $D=1
M5 15 15 4 4 nmos_a L=2.4e-07 W=1.2e-06 AD=7.2e-13 AS=4.8e-13 PD=1.8e-06 PS=9e-07 w_cont=6e-07 nfing=1 source_num=2 $X=-132740 $Y=-144820 $D=1
M6 16 16 17 17 nmos_a L=2.4e-07 W=1.2e-06 AD=7.2e-13 AS=4.8e-13 PD=1.8e-06 PS=9e-07 w_cont=6e-07 nfing=1 source_num=2 $X=-112940 $Y=-144820 $D=1
M7 18 18 4 4 nmos_a L=2.4e-07 W=1.2e-06 AD=7.2e-13 AS=4.8e-13 PD=1.8e-06 PS=9e-07 w_cont=6e-07 nfing=1 source_num=2 $X=-107540 $Y=-144820 $D=1
M8 19 19 20 20 nmos_a L=2.4e-07 W=1.2e-06 AD=7.2e-13 AS=4.8e-13 PD=1.8e-06 PS=9e-07 w_cont=6e-07 nfing=1 source_num=2 $X=-87740 $Y=-144820 $D=1
M9 21 21 4 4 nmos_a L=2.4e-07 W=1.2e-06 AD=7.2e-13 AS=4.8e-13 PD=1.8e-06 PS=9e-07 w_cont=6e-07 nfing=1 source_num=2 $X=-82340 $Y=-144820 $D=1
X10 5 7 7 pmos_a_CDNS_5887047866540 $T=-189240 -143960 1 270 $X=-191440 $Y=-145400
X11 8 9 9 pmos_a_CDNS_5887047866540 $T=-183840 -143960 1 270 $X=-186040 $Y=-145400
X12 5 3 5 pmos_a_CDNS_5887047866540 $T=-178300 -145440 0 90 $X=-180500 $Y=-145440
X13 5 10 10 pmos_a_CDNS_5887047866540 $T=-164040 -143960 1 270 $X=-166240 $Y=-145400
X14 11 12 12 pmos_a_CDNS_5887047866540 $T=-158640 -143960 1 270 $X=-160840 $Y=-145400
X15 5 3 5 pmos_a_CDNS_5887047866540 $T=-153100 -145440 0 90 $X=-155300 $Y=-145440
X16 5 13 13 pmos_a_CDNS_5887047866540 $T=-138840 -143960 1 270 $X=-141040 $Y=-145400
X17 14 15 15 pmos_a_CDNS_5887047866540 $T=-133440 -143960 1 270 $X=-135640 $Y=-145400
X18 5 3 5 pmos_a_CDNS_5887047866540 $T=-127900 -145440 0 90 $X=-130100 $Y=-145440
X19 5 16 16 pmos_a_CDNS_5887047866540 $T=-113640 -143960 1 270 $X=-115840 $Y=-145400
X20 17 18 18 pmos_a_CDNS_5887047866540 $T=-108240 -143960 1 270 $X=-110440 $Y=-145400
X21 5 3 5 pmos_a_CDNS_5887047866540 $T=-102700 -145440 0 90 $X=-104900 $Y=-145440
X22 5 19 19 pmos_a_CDNS_5887047866540 $T=-88440 -143960 1 270 $X=-90640 $Y=-145400
X23 20 21 21 pmos_a_CDNS_5887047866540 $T=-83040 -143960 1 270 $X=-85240 $Y=-145400
X34 3 2 5 nmos_a_CDNS_5887047866547 $T=-177720 -143960 0 270 $X=-177720 $Y=-145400
X35 3 2 5 nmos_a_CDNS_5887047866547 $T=-152520 -143960 0 270 $X=-152520 $Y=-145400
X36 3 2 5 nmos_a_CDNS_5887047866547 $T=-127320 -143960 0 270 $X=-127320 $Y=-145400
X37 3 2 5 nmos_a_CDNS_5887047866547 $T=-102120 -143960 0 270 $X=-102120 $Y=-145400
.ENDS
***************************************
.SUBCKT pmos_a_CDNS_5887047866560
** N=3 EP=0 IP=0 FDC=0
*.SEEDPROM
.ENDS
***************************************
.SUBCKT nmos_a_CDNS_5887047866554
** N=3 EP=0 IP=0 FDC=0
*.SEEDPROM
.ENDS
***************************************
.SUBCKT Cell_Usub Low nmos pmos High
** N=4 EP=4 IP=0 FDC=4
*.SEEDPROM
M0 nmos Low Low Low nmos_a L=3.8e-07 W=4.8e-07 AD=4.24e-13 AS=1.92e-13 PD=1.06e-06 PS=5.3e-07 w_cont=5.8e-07 nfing=1 source_num=2 $X=1280 $Y=2220 $D=1
M1 nmos Low Low Low nmos_a L=3.8e-07 W=4.8e-07 AD=4.24e-13 AS=1.92e-13 PD=1.06e-06 PS=5.3e-07 w_cont=5.8e-07 nfing=1 source_num=2 $X=3700 $Y=2220 $D=1
M2 pmos High High High pmos_h L=2.4e-07 W=6.6e-07 AD=2.64e-13 AS=2.64e-13 PD=1.46e-06 PS=1.46e-06 m=1 $X=1860 $Y=760 $D=6
M3 pmos High High High pmos_h L=2.4e-07 W=6.6e-07 AD=2.64e-13 AS=2.64e-13 PD=1.46e-06 PS=1.46e-06 m=1 $X=3520 $Y=760 $D=6
.ENDS
***************************************
.SUBCKT ICV_149 1 2 3 4
** N=4 EP=4 IP=8 FDC=10
*.SEEDPROM
M0 1 4 4 4 pmos_a L=2.4e-07 W=1e-06 AD=5.928e-13 AS=1.61e-13 PD=1.6e-06 PS=8e-07 w_cont=6e-07 nfing=1 mmm=1 $X=5540 $Y=360 $D=5
M1 1 4 4 4 pmos_a L=2.4e-07 W=1e-06 AD=5.928e-13 AS=1.61e-13 PD=1.6e-06 PS=8e-07 w_cont=6e-07 nfing=1 mmm=1 $X=6300 $Y=360 $D=5
X2 3 2 1 4 Cell_Usub $T=0 0 0 0 $X=-360 $Y=-340
X3 3 2 1 4 Cell_Usub $T=6040 0 0 0 $X=5680 $Y=-340
.ENDS
***************************************
.SUBCKT ICV_150 1 2 3 4
** N=4 EP=4 IP=8 FDC=23
*.SEEDPROM
M0 1 4 4 4 pmos_a L=2.4e-07 W=1e-06 AD=5.928e-13 AS=1.61e-13 PD=1.6e-06 PS=8e-07 w_cont=6e-07 nfing=1 mmm=1 $X=260 $Y=360 $D=5
M1 1 4 4 4 pmos_a L=2.4e-07 W=1e-06 AD=5.928e-13 AS=1.61e-13 PD=1.6e-06 PS=8e-07 w_cont=6e-07 nfing=1 mmm=1 $X=11580 $Y=360 $D=5
M2 1 4 4 4 pmos_a L=2.4e-07 W=1e-06 AD=5.928e-13 AS=1.61e-13 PD=1.6e-06 PS=8e-07 w_cont=6e-07 nfing=1 mmm=1 $X=12340 $Y=360 $D=5
X3 1 2 3 4 ICV_149 $T=0 0 0 0 $X=-360 $Y=-340
X4 1 2 3 4 ICV_149 $T=12080 0 0 0 $X=11720 $Y=-340
.ENDS
***************************************
.SUBCKT ICV_151 1 2 3 4 5 6 7 8 9 10 11 12 13 14 15 16 17 18
** N=22 EP=18 IP=224 FDC=559
*.SEEDPROM
M0 1 4 1 1 nmos_a L=2e-06 W=5.5e-06 AD=8.30487e-13 AS=2.2e-12 PD=1.59709e-06 PS=1.59709e-06 w_cont=6e-07 nfing=1 source_num=2 $X=-213980 $Y=275380 $D=1
M1 1 4 1 1 nmos_a L=2e-06 W=5.5e-06 AD=8.30487e-13 AS=1.43e-12 PD=1.59709e-06 PS=1.59709e-06 w_cont=6e-07 nfing=1 source_num=2 $X=-211460 $Y=275380 $D=1
M2 1 4 1 1 nmos_a L=2e-06 W=5.5e-06 AD=8.30487e-13 AS=1.43e-12 PD=1.59709e-06 PS=1.59709e-06 w_cont=6e-07 nfing=1 source_num=2 $X=-208940 $Y=275380 $D=1
M3 1 4 1 1 nmos_a L=2e-06 W=5.5e-06 AD=8.30487e-13 AS=1.43e-12 PD=1.59709e-06 PS=1.59709e-06 w_cont=6e-07 nfing=1 source_num=2 $X=-206420 $Y=275380 $D=1
M4 1 4 1 1 nmos_a L=2e-06 W=5.5e-06 AD=8.30487e-13 AS=1.43e-12 PD=1.59709e-06 PS=1.59709e-06 w_cont=6e-07 nfing=1 source_num=2 $X=-203900 $Y=275380 $D=1
M5 11 6 1 1 nmos_a L=2.4e-07 W=1.2e-06 AD=4.68e-13 AS=4.8e-13 PD=9e-07 PS=9e-07 w_cont=6e-07 nfing=1 source_num=2 $X=-203700 $Y=271520 $D=1
M6 11 6 1 1 nmos_a L=2.4e-07 W=1.2e-06 AD=4.68e-13 AS=4.8e-13 PD=9e-07 PS=9e-07 w_cont=6e-07 nfing=1 source_num=2 $X=-202940 $Y=271520 $D=1
M7 1 4 1 1 nmos_a L=2e-06 W=5.5e-06 AD=8.30487e-13 AS=1.43e-12 PD=1.59709e-06 PS=1.59709e-06 w_cont=6e-07 nfing=1 source_num=2 $X=-201380 $Y=275380 $D=1
M8 14 5 21 21 nmos_a L=4.8e-07 W=4.8e-07 AD=7.128e-13 AS=2.304e-13 PD=1.08e-06 PS=5.4e-07 w_cont=6e-07 nfing=1 source_num=2 $X=-200840 $Y=270140 $D=1
M9 1 4 1 1 nmos_a L=2e-06 W=5.5e-06 AD=8.30487e-13 AS=1.43e-12 PD=1.59709e-06 PS=1.59709e-06 w_cont=6e-07 nfing=1 source_num=2 $X=-198860 $Y=275380 $D=1
M10 14 13 1 1 nmos_a L=4.8e-07 W=4.8e-07 AD=4.32e-13 AS=2.496e-13 PD=1.08e-06 PS=5.4e-07 w_cont=6e-07 nfing=1 source_num=2 $X=-198540 $Y=272160 $D=1
M11 15 14 1 1 nmos_a L=2.4e-07 W=4.8e-07 AD=4.32e-13 AS=2.496e-13 PD=1.08e-06 PS=5.4e-07 w_cont=6e-07 nfing=1 source_num=2 $X=-197540 $Y=272160 $D=1
M12 6 15 16 16 nmos_a L=2.4e-07 W=4.8e-07 AD=4.32e-13 AS=1.92e-13 PD=1.08e-06 PS=5.4e-07 w_cont=6e-07 nfing=1 source_num=2 $X=-195880 $Y=272160 $D=1
M13 10 3 20 20 nmos_a L=3e-07 W=1.2e-06 AD=7.2e-13 AS=6.24e-13 PD=1.8e-06 PS=9e-07 w_cont=6e-07 nfing=1 source_num=2 $X=-213020 $Y=269000 $D=1
M14 5 9 20 20 nmos_a L=3e-07 W=1.2e-06 AD=7.2e-13 AS=6.24e-13 PD=1.8e-06 PS=9e-07 w_cont=6e-07 nfing=1 source_num=2 $X=-212200 $Y=269000 $D=1
M15 20 4 1 1 nmos_a L=3e-07 W=1.2e-06 AD=7.2e-13 AS=3.12e-13 PD=1.8e-06 PS=9e-07 w_cont=6e-07 nfing=1 source_num=2 $X=-212240 $Y=272640 $D=1
M16 4 4 1 1 nmos_a L=3e-07 W=1.2e-06 AD=7.2e-13 AS=3.12e-13 PD=1.8e-06 PS=9e-07 w_cont=6e-07 nfing=1 source_num=2 $X=-211420 $Y=272640 $D=1
M17 10 3 20 20 nmos_a L=3e-07 W=1.2e-06 AD=7.2e-13 AS=6.24e-13 PD=1.8e-06 PS=9e-07 w_cont=6e-07 nfing=1 source_num=2 $X=-210700 $Y=269000 $D=1
M18 5 9 20 20 nmos_a L=3e-07 W=1.2e-06 AD=7.2e-13 AS=6.24e-13 PD=1.8e-06 PS=9e-07 w_cont=6e-07 nfing=1 source_num=2 $X=-209880 $Y=269000 $D=1
M19 20 4 1 1 nmos_a L=3e-07 W=1.2e-06 AD=7.2e-13 AS=4.8e-13 PD=1.8e-06 PS=9e-07 w_cont=6e-07 nfing=1 source_num=2 $X=-209920 $Y=272640 $D=1
M20 10 3 20 20 nmos_a L=3e-07 W=1.2e-06 AD=7.2e-13 AS=6.24e-13 PD=1.8e-06 PS=9e-07 w_cont=6e-07 nfing=1 source_num=2 $X=-208380 $Y=269000 $D=1
M21 20 4 1 1 nmos_a L=3e-07 W=1.2e-06 AD=7.2e-13 AS=3.12e-13 PD=1.8e-06 PS=9e-07 w_cont=6e-07 nfing=1 source_num=2 $X=-208380 $Y=272640 $D=1
M22 5 9 20 20 nmos_a L=3e-07 W=1.2e-06 AD=7.2e-13 AS=6.24e-13 PD=1.8e-06 PS=9e-07 w_cont=6e-07 nfing=1 source_num=2 $X=-207560 $Y=269000 $D=1
M23 4 4 1 1 nmos_a L=3e-07 W=1.2e-06 AD=7.2e-13 AS=3.12e-13 PD=1.8e-06 PS=9e-07 w_cont=6e-07 nfing=1 source_num=2 $X=-207560 $Y=272640 $D=1
M24 10 3 20 20 nmos_a L=3e-07 W=1.2e-06 AD=7.2e-13 AS=6.24e-13 PD=1.8e-06 PS=9e-07 w_cont=6e-07 nfing=1 source_num=2 $X=-206060 $Y=269000 $D=1
M25 20 4 1 1 nmos_a L=3e-07 W=1.2e-06 AD=7.2e-13 AS=4.8e-13 PD=1.8e-06 PS=9e-07 w_cont=6e-07 nfing=1 source_num=2 $X=-206060 $Y=272640 $D=1
M26 5 9 20 20 nmos_a L=3e-07 W=1.2e-06 AD=7.2e-13 AS=6.24e-13 PD=1.8e-06 PS=9e-07 w_cont=6e-07 nfing=1 source_num=2 $X=-205240 $Y=269000 $D=1
M27 21 4 1 1 nmos_a L=3e-07 W=1.2e-06 AD=7.2e-13 AS=4.8e-13 PD=1.8e-06 PS=9e-07 w_cont=6e-07 nfing=1 source_num=2 $X=-201500 $Y=272200 $D=1
M28 12 4 13 13 nmos_a L=3e-07 W=1.2e-06 AD=7.2e-13 AS=4.8e-13 PD=1.8e-06 PS=9e-07 w_cont=6e-07 nfing=1 source_num=2 $X=-200040 $Y=272200 $D=1
M29 9 7 1 1 nmos_a L=3e-07 W=4.8e-07 AD=2.808e-13 AS=1.92e-13 PD=5.4e-07 PS=5.4e-07 w_cont=6e-07 nfing=1 source_num=2 $X=-223460 $Y=268220 $D=1
M30 9 7 1 1 nmos_a L=3e-07 W=4.8e-07 AD=2.808e-13 AS=1.248e-13 PD=5.4e-07 PS=5.4e-07 w_cont=6e-07 nfing=1 source_num=2 $X=-222640 $Y=268220 $D=1
M31 9 7 1 1 nmos_a L=3e-07 W=4.8e-07 AD=2.808e-13 AS=1.248e-13 PD=5.4e-07 PS=5.4e-07 w_cont=6e-07 nfing=1 source_num=2 $X=-221820 $Y=268220 $D=1
M32 9 7 1 1 nmos_a L=3e-07 W=4.8e-07 AD=2.808e-13 AS=1.248e-13 PD=5.4e-07 PS=5.4e-07 w_cont=6e-07 nfing=1 source_num=2 $X=-221000 $Y=268220 $D=1
M33 9 7 1 1 nmos_a L=3e-07 W=4.8e-07 AD=2.808e-13 AS=1.248e-13 PD=5.4e-07 PS=5.4e-07 w_cont=6e-07 nfing=1 source_num=2 $X=-220180 $Y=268220 $D=1
M34 9 7 1 1 nmos_a L=3e-07 W=4.8e-07 AD=2.808e-13 AS=1.248e-13 PD=5.4e-07 PS=5.4e-07 w_cont=6e-07 nfing=1 source_num=2 $X=-219360 $Y=268220 $D=1
M35 9 7 1 1 nmos_a L=3e-07 W=4.8e-07 AD=2.808e-13 AS=1.248e-13 PD=5.4e-07 PS=5.4e-07 w_cont=6e-07 nfing=1 source_num=2 $X=-218540 $Y=268220 $D=1
M36 9 7 1 1 nmos_a L=3e-07 W=4.8e-07 AD=2.808e-13 AS=1.248e-13 PD=5.4e-07 PS=5.4e-07 w_cont=6e-07 nfing=1 source_num=2 $X=-217720 $Y=268220 $D=1
M37 9 7 1 1 nmos_a L=3e-07 W=4.8e-07 AD=2.808e-13 AS=1.248e-13 PD=5.4e-07 PS=5.4e-07 w_cont=6e-07 nfing=1 source_num=2 $X=-216900 $Y=268220 $D=1
M38 9 7 1 1 nmos_a L=3e-07 W=4.8e-07 AD=2.808e-13 AS=1.92e-13 PD=5.4e-07 PS=5.4e-07 w_cont=6e-07 nfing=1 source_num=2 $X=-216080 $Y=268220 $D=1
M39 22 12 2 2 pmos_a L=2.4e-07 W=4.8e-07 AD=4.32e-13 AS=1.224e-13 PD=1.08e-06 PS=5.4e-07 w_cont=6e-07 nfing=1 mmm=1 $X=-199120 $Y=269000 $D=5
M40 14 5 22 22 pmos_a L=2.4e-07 W=4.8e-07 AD=4.32e-13 AS=1.584e-13 PD=1.08e-06 PS=5.4e-07 w_cont=6e-07 nfing=1 mmm=1 $X=-199120 $Y=270380 $D=5
M41 14 15 22 22 pmos_a L=2.4e-07 W=4.8e-07 AD=4.32e-13 AS=1.584e-13 PD=1.08e-06 PS=5.4e-07 w_cont=6e-07 nfing=1 mmm=1 $X=-199120 $Y=271140 $D=5
M42 9 8 2 2 pmos_a L=3e-07 W=4.8e-07 AD=2.808e-13 AS=1.224e-13 PD=5.4e-07 PS=5.4e-07 w_cont=6e-07 nfing=1 mmm=1 $X=-223460 $Y=270500 $D=5
M43 9 8 2 2 pmos_a L=3e-07 W=4.8e-07 AD=2.808e-13 AS=1.224e-13 PD=5.4e-07 PS=5.4e-07 w_cont=6e-07 nfing=1 mmm=1 $X=-223460 $Y=271980 $D=5
M44 9 8 2 2 pmos_a L=3e-07 W=4.8e-07 AD=2.808e-13 AS=1.224e-13 PD=5.4e-07 PS=5.4e-07 w_cont=6e-07 nfing=1 mmm=1 $X=-223460 $Y=273460 $D=5
M45 9 8 2 2 pmos_a L=3e-07 W=4.8e-07 AD=2.808e-13 AS=1.584e-13 PD=5.4e-07 PS=5.4e-07 w_cont=6e-07 nfing=1 mmm=1 $X=-222640 $Y=270500 $D=5
M46 9 8 2 2 pmos_a L=3e-07 W=4.8e-07 AD=2.808e-13 AS=1.584e-13 PD=5.4e-07 PS=5.4e-07 w_cont=6e-07 nfing=1 mmm=1 $X=-222640 $Y=271980 $D=5
M47 9 8 2 2 pmos_a L=3e-07 W=4.8e-07 AD=2.808e-13 AS=1.584e-13 PD=5.4e-07 PS=5.4e-07 w_cont=6e-07 nfing=1 mmm=1 $X=-222640 $Y=273460 $D=5
M48 9 8 2 2 pmos_a L=3e-07 W=4.8e-07 AD=2.808e-13 AS=1.584e-13 PD=5.4e-07 PS=5.4e-07 w_cont=6e-07 nfing=1 mmm=1 $X=-221820 $Y=270500 $D=5
M49 9 8 2 2 pmos_a L=3e-07 W=4.8e-07 AD=2.808e-13 AS=1.584e-13 PD=5.4e-07 PS=5.4e-07 w_cont=6e-07 nfing=1 mmm=1 $X=-221820 $Y=271980 $D=5
M50 8 8 2 2 pmos_a L=3e-07 W=4.8e-07 AD=2.808e-13 AS=1.584e-13 PD=5.4e-07 PS=5.4e-07 w_cont=6e-07 nfing=1 mmm=1 $X=-221820 $Y=273460 $D=5
M51 9 8 2 2 pmos_a L=3e-07 W=4.8e-07 AD=2.808e-13 AS=1.584e-13 PD=5.4e-07 PS=5.4e-07 w_cont=6e-07 nfing=1 mmm=1 $X=-221000 $Y=270500 $D=5
M52 9 8 2 2 pmos_a L=3e-07 W=4.8e-07 AD=2.808e-13 AS=1.584e-13 PD=5.4e-07 PS=5.4e-07 w_cont=6e-07 nfing=1 mmm=1 $X=-221000 $Y=271980 $D=5
M53 8 8 2 2 pmos_a L=3e-07 W=4.8e-07 AD=2.808e-13 AS=1.584e-13 PD=5.4e-07 PS=5.4e-07 w_cont=6e-07 nfing=1 mmm=1 $X=-221000 $Y=273460 $D=5
M54 9 8 2 2 pmos_a L=3e-07 W=4.8e-07 AD=2.808e-13 AS=1.584e-13 PD=5.4e-07 PS=5.4e-07 w_cont=6e-07 nfing=1 mmm=1 $X=-220180 $Y=270500 $D=5
M55 9 8 2 2 pmos_a L=3e-07 W=4.8e-07 AD=2.808e-13 AS=1.584e-13 PD=5.4e-07 PS=5.4e-07 w_cont=6e-07 nfing=1 mmm=1 $X=-220180 $Y=271980 $D=5
M56 9 8 2 2 pmos_a L=3e-07 W=4.8e-07 AD=2.808e-13 AS=1.584e-13 PD=5.4e-07 PS=5.4e-07 w_cont=6e-07 nfing=1 mmm=1 $X=-220180 $Y=273460 $D=5
M57 9 8 2 2 pmos_a L=3e-07 W=4.8e-07 AD=2.808e-13 AS=1.584e-13 PD=5.4e-07 PS=5.4e-07 w_cont=6e-07 nfing=1 mmm=1 $X=-219360 $Y=270500 $D=5
M58 9 8 2 2 pmos_a L=3e-07 W=4.8e-07 AD=2.808e-13 AS=1.584e-13 PD=5.4e-07 PS=5.4e-07 w_cont=6e-07 nfing=1 mmm=1 $X=-219360 $Y=271980 $D=5
M59 9 8 2 2 pmos_a L=3e-07 W=4.8e-07 AD=2.808e-13 AS=1.584e-13 PD=5.4e-07 PS=5.4e-07 w_cont=6e-07 nfing=1 mmm=1 $X=-219360 $Y=273460 $D=5
M60 9 8 2 2 pmos_a L=3e-07 W=4.8e-07 AD=2.808e-13 AS=1.584e-13 PD=5.4e-07 PS=5.4e-07 w_cont=6e-07 nfing=1 mmm=1 $X=-218540 $Y=270500 $D=5
M61 9 8 2 2 pmos_a L=3e-07 W=4.8e-07 AD=2.808e-13 AS=1.584e-13 PD=5.4e-07 PS=5.4e-07 w_cont=6e-07 nfing=1 mmm=1 $X=-218540 $Y=271980 $D=5
M62 8 8 2 2 pmos_a L=3e-07 W=4.8e-07 AD=2.808e-13 AS=1.584e-13 PD=5.4e-07 PS=5.4e-07 w_cont=6e-07 nfing=1 mmm=1 $X=-218540 $Y=273460 $D=5
M63 9 8 2 2 pmos_a L=3e-07 W=4.8e-07 AD=2.808e-13 AS=1.584e-13 PD=5.4e-07 PS=5.4e-07 w_cont=6e-07 nfing=1 mmm=1 $X=-217720 $Y=270500 $D=5
M64 9 8 2 2 pmos_a L=3e-07 W=4.8e-07 AD=2.808e-13 AS=1.584e-13 PD=5.4e-07 PS=5.4e-07 w_cont=6e-07 nfing=1 mmm=1 $X=-217720 $Y=271980 $D=5
M65 8 8 2 2 pmos_a L=3e-07 W=4.8e-07 AD=2.808e-13 AS=1.584e-13 PD=5.4e-07 PS=5.4e-07 w_cont=6e-07 nfing=1 mmm=1 $X=-217720 $Y=273460 $D=5
M66 9 8 2 2 pmos_a L=3e-07 W=4.8e-07 AD=2.808e-13 AS=1.584e-13 PD=5.4e-07 PS=5.4e-07 w_cont=6e-07 nfing=1 mmm=1 $X=-216900 $Y=270500 $D=5
M67 9 8 2 2 pmos_a L=3e-07 W=4.8e-07 AD=2.808e-13 AS=1.584e-13 PD=5.4e-07 PS=5.4e-07 w_cont=6e-07 nfing=1 mmm=1 $X=-216900 $Y=271980 $D=5
M68 9 8 2 2 pmos_a L=3e-07 W=4.8e-07 AD=2.808e-13 AS=1.584e-13 PD=5.4e-07 PS=5.4e-07 w_cont=6e-07 nfing=1 mmm=1 $X=-216900 $Y=273460 $D=5
M69 9 8 2 2 pmos_a L=3e-07 W=4.8e-07 AD=2.808e-13 AS=1.224e-13 PD=5.4e-07 PS=5.4e-07 w_cont=6e-07 nfing=1 mmm=1 $X=-216080 $Y=270500 $D=5
M70 9 8 2 2 pmos_a L=3e-07 W=4.8e-07 AD=2.808e-13 AS=1.224e-13 PD=5.4e-07 PS=5.4e-07 w_cont=6e-07 nfing=1 mmm=1 $X=-216080 $Y=271980 $D=5
M71 9 8 2 2 pmos_a L=3e-07 W=4.8e-07 AD=2.808e-13 AS=1.224e-13 PD=5.4e-07 PS=5.4e-07 w_cont=6e-07 nfing=1 mmm=1 $X=-216080 $Y=273460 $D=5
M72 7 18 18 18 pmos_a L=2.4e-07 W=1e-06 AD=5.928e-13 AS=1.61e-13 PD=1.6e-06 PS=8e-07 w_cont=6e-07 nfing=1 mmm=1 $X=-372180 $Y=269800 $D=5
M73 7 18 18 18 pmos_a L=2.4e-07 W=1e-06 AD=5.928e-13 AS=1.61e-13 PD=1.6e-06 PS=8e-07 w_cont=6e-07 nfing=1 mmm=1 $X=-372180 $Y=272120 $D=5
M74 7 18 18 18 pmos_a L=2.4e-07 W=1e-06 AD=5.928e-13 AS=1.61e-13 PD=1.6e-06 PS=8e-07 w_cont=6e-07 nfing=1 mmm=1 $X=-348020 $Y=269800 $D=5
M75 7 18 18 18 pmos_a L=2.4e-07 W=1e-06 AD=5.928e-13 AS=1.61e-13 PD=1.6e-06 PS=8e-07 w_cont=6e-07 nfing=1 mmm=1 $X=-348020 $Y=272120 $D=5
M76 7 18 18 18 pmos_a L=2.4e-07 W=1e-06 AD=5.928e-13 AS=1.61e-13 PD=1.6e-06 PS=8e-07 w_cont=6e-07 nfing=1 mmm=1 $X=-323860 $Y=269800 $D=5
M77 7 18 18 18 pmos_a L=2.4e-07 W=1e-06 AD=5.928e-13 AS=1.61e-13 PD=1.6e-06 PS=8e-07 w_cont=6e-07 nfing=1 mmm=1 $X=-323860 $Y=272120 $D=5
M78 7 18 18 18 pmos_a L=2.4e-07 W=1e-06 AD=5.928e-13 AS=1.61e-13 PD=1.6e-06 PS=8e-07 w_cont=6e-07 nfing=1 mmm=1 $X=-299700 $Y=269800 $D=5
M79 7 18 18 18 pmos_a L=2.4e-07 W=1e-06 AD=5.928e-13 AS=1.61e-13 PD=1.6e-06 PS=8e-07 w_cont=6e-07 nfing=1 mmm=1 $X=-299700 $Y=272120 $D=5
M80 7 18 18 18 pmos_a L=2.4e-07 W=1e-06 AD=5.928e-13 AS=1.61e-13 PD=1.6e-06 PS=8e-07 w_cont=6e-07 nfing=1 mmm=1 $X=-275540 $Y=269800 $D=5
M81 7 18 18 18 pmos_a L=2.4e-07 W=1e-06 AD=5.928e-13 AS=1.61e-13 PD=1.6e-06 PS=8e-07 w_cont=6e-07 nfing=1 mmm=1 $X=-275540 $Y=272120 $D=5
M82 7 18 18 18 pmos_a L=2.4e-07 W=1e-06 AD=5.928e-13 AS=1.61e-13 PD=1.6e-06 PS=8e-07 w_cont=6e-07 nfing=1 mmm=1 $X=-251380 $Y=269800 $D=5
M83 7 18 18 18 pmos_a L=2.4e-07 W=1e-06 AD=5.928e-13 AS=1.61e-13 PD=1.6e-06 PS=8e-07 w_cont=6e-07 nfing=1 mmm=1 $X=-251380 $Y=272120 $D=5
M84 7 18 18 18 pmos_a L=2.4e-07 W=1e-06 AD=5.928e-13 AS=1.25e-13 PD=1.6e-06 PS=8e-07 w_cont=6e-07 nfing=1 mmm=1 $X=-227220 $Y=269800 $D=5
M85 7 18 18 18 pmos_a L=2.4e-07 W=1e-06 AD=5.928e-13 AS=1.25e-13 PD=1.6e-06 PS=8e-07 w_cont=6e-07 nfing=1 mmm=1 $X=-227220 $Y=272120 $D=5
M86 1 2 1 cpoly_p w=3.8e-06 l=2e-06 c=5.2038e-14 as=2.31158e-13 ad=7.488e-13 ps=1.44e-06 pd=1.11673e-06 sim_w=2.88e-06 m_per_maxw=1.31944 numb_sub_cont=3 nfing=1 $X=-396100 $Y=276580 $D=21
M87 1 2 1 cpoly_p w=3.8e-06 l=2e-06 c=5.2038e-14 as=2.31158e-13 ad=7.488e-13 ps=1.44e-06 pd=1.11673e-06 sim_w=2.88e-06 m_per_maxw=1.31944 numb_sub_cont=3 nfing=1 $X=-393580 $Y=276580 $D=21
M88 1 2 1 cpoly_p w=3.8e-06 l=2e-06 c=5.2038e-14 as=2.31158e-13 ad=7.488e-13 ps=1.44e-06 pd=1.11673e-06 sim_w=2.88e-06 m_per_maxw=1.31944 numb_sub_cont=3 nfing=1 $X=-391060 $Y=276580 $D=21
M89 1 2 1 cpoly_p w=3.8e-06 l=2e-06 c=5.2038e-14 as=2.31158e-13 ad=7.488e-13 ps=1.44e-06 pd=1.11673e-06 sim_w=2.88e-06 m_per_maxw=1.31944 numb_sub_cont=3 nfing=1 $X=-388540 $Y=276580 $D=21
M90 1 2 1 cpoly_p w=3.8e-06 l=2e-06 c=5.2038e-14 as=2.31158e-13 ad=7.488e-13 ps=1.44e-06 pd=1.11673e-06 sim_w=2.88e-06 m_per_maxw=1.31944 numb_sub_cont=3 nfing=1 $X=-386020 $Y=276580 $D=21
M91 1 2 1 cpoly_p w=3.8e-06 l=2e-06 c=5.2038e-14 as=2.31158e-13 ad=7.488e-13 ps=1.44e-06 pd=1.11673e-06 sim_w=2.88e-06 m_per_maxw=1.31944 numb_sub_cont=3 nfing=1 $X=-383500 $Y=276580 $D=21
M92 1 2 1 cpoly_p w=3.8e-06 l=2e-06 c=5.2038e-14 as=2.31158e-13 ad=7.488e-13 ps=1.44e-06 pd=1.11673e-06 sim_w=2.88e-06 m_per_maxw=1.31944 numb_sub_cont=3 nfing=1 $X=-380980 $Y=276580 $D=21
M93 1 2 1 cpoly_p w=3.8e-06 l=2e-06 c=5.2038e-14 as=2.31158e-13 ad=7.488e-13 ps=1.44e-06 pd=1.11673e-06 sim_w=2.88e-06 m_per_maxw=1.31944 numb_sub_cont=3 nfing=1 $X=-378460 $Y=276580 $D=21
M94 1 2 1 cpoly_p w=3.8e-06 l=2e-06 c=5.2038e-14 as=2.31158e-13 ad=7.488e-13 ps=1.44e-06 pd=1.11673e-06 sim_w=2.88e-06 m_per_maxw=1.31944 numb_sub_cont=3 nfing=1 $X=-375940 $Y=276580 $D=21
M95 1 2 1 cpoly_p w=3.8e-06 l=2e-06 c=5.2038e-14 as=2.31158e-13 ad=7.488e-13 ps=1.44e-06 pd=1.11673e-06 sim_w=2.88e-06 m_per_maxw=1.31944 numb_sub_cont=3 nfing=1 $X=-373420 $Y=276580 $D=21
M96 1 2 1 cpoly_p w=3.8e-06 l=2e-06 c=5.2038e-14 as=2.31158e-13 ad=7.488e-13 ps=1.44e-06 pd=1.11673e-06 sim_w=2.88e-06 m_per_maxw=1.31944 numb_sub_cont=3 nfing=1 $X=-370900 $Y=276580 $D=21
M97 1 2 1 cpoly_p w=3.8e-06 l=2e-06 c=5.2038e-14 as=2.31158e-13 ad=7.488e-13 ps=1.44e-06 pd=1.11673e-06 sim_w=2.88e-06 m_per_maxw=1.31944 numb_sub_cont=3 nfing=1 $X=-368380 $Y=276580 $D=21
M98 1 2 1 cpoly_p w=3.8e-06 l=2e-06 c=5.2038e-14 as=2.31158e-13 ad=7.488e-13 ps=1.44e-06 pd=1.11673e-06 sim_w=2.88e-06 m_per_maxw=1.31944 numb_sub_cont=3 nfing=1 $X=-365860 $Y=276580 $D=21
M99 1 2 1 cpoly_p w=3.8e-06 l=2e-06 c=5.2038e-14 as=2.31158e-13 ad=7.488e-13 ps=1.44e-06 pd=1.11673e-06 sim_w=2.88e-06 m_per_maxw=1.31944 numb_sub_cont=3 nfing=1 $X=-363340 $Y=276580 $D=21
M100 1 2 1 cpoly_p w=3.8e-06 l=2e-06 c=5.2038e-14 as=2.31158e-13 ad=7.488e-13 ps=1.44e-06 pd=1.11673e-06 sim_w=2.88e-06 m_per_maxw=1.31944 numb_sub_cont=3 nfing=1 $X=-360820 $Y=276580 $D=21
M101 1 2 1 cpoly_p w=3.8e-06 l=2e-06 c=5.2038e-14 as=2.31158e-13 ad=7.488e-13 ps=1.44e-06 pd=1.11673e-06 sim_w=2.88e-06 m_per_maxw=1.31944 numb_sub_cont=3 nfing=1 $X=-358300 $Y=276580 $D=21
M102 1 2 1 cpoly_p w=3.8e-06 l=2e-06 c=5.2038e-14 as=2.31158e-13 ad=7.488e-13 ps=1.44e-06 pd=1.11673e-06 sim_w=2.88e-06 m_per_maxw=1.31944 numb_sub_cont=3 nfing=1 $X=-355780 $Y=276580 $D=21
M103 1 2 1 cpoly_p w=3.8e-06 l=2e-06 c=5.2038e-14 as=2.31158e-13 ad=7.488e-13 ps=1.44e-06 pd=1.11673e-06 sim_w=2.88e-06 m_per_maxw=1.31944 numb_sub_cont=3 nfing=1 $X=-353260 $Y=276580 $D=21
M104 1 2 1 cpoly_p w=3.8e-06 l=2e-06 c=5.2038e-14 as=2.31158e-13 ad=7.488e-13 ps=1.44e-06 pd=1.11673e-06 sim_w=2.88e-06 m_per_maxw=1.31944 numb_sub_cont=3 nfing=1 $X=-350740 $Y=276580 $D=21
M105 1 2 1 cpoly_p w=3.8e-06 l=2e-06 c=5.2038e-14 as=2.31158e-13 ad=7.488e-13 ps=1.44e-06 pd=1.11673e-06 sim_w=2.88e-06 m_per_maxw=1.31944 numb_sub_cont=3 nfing=1 $X=-348220 $Y=276580 $D=21
M106 1 2 1 cpoly_p w=3.8e-06 l=2e-06 c=5.2038e-14 as=2.31158e-13 ad=7.488e-13 ps=1.44e-06 pd=1.11673e-06 sim_w=2.88e-06 m_per_maxw=1.31944 numb_sub_cont=3 nfing=1 $X=-345700 $Y=276580 $D=21
M107 1 2 1 cpoly_p w=3.8e-06 l=2e-06 c=5.2038e-14 as=2.31158e-13 ad=7.488e-13 ps=1.44e-06 pd=1.11673e-06 sim_w=2.88e-06 m_per_maxw=1.31944 numb_sub_cont=3 nfing=1 $X=-343180 $Y=276580 $D=21
M108 1 2 1 cpoly_p w=3.8e-06 l=2e-06 c=5.2038e-14 as=2.31158e-13 ad=7.488e-13 ps=1.44e-06 pd=1.11673e-06 sim_w=2.88e-06 m_per_maxw=1.31944 numb_sub_cont=3 nfing=1 $X=-340660 $Y=276580 $D=21
M109 1 2 1 cpoly_p w=3.8e-06 l=2e-06 c=5.2038e-14 as=2.31158e-13 ad=7.488e-13 ps=1.44e-06 pd=1.11673e-06 sim_w=2.88e-06 m_per_maxw=1.31944 numb_sub_cont=3 nfing=1 $X=-338140 $Y=276580 $D=21
M110 1 2 1 cpoly_p w=3.8e-06 l=2e-06 c=5.2038e-14 as=2.31158e-13 ad=7.488e-13 ps=1.44e-06 pd=1.11673e-06 sim_w=2.88e-06 m_per_maxw=1.31944 numb_sub_cont=3 nfing=1 $X=-335620 $Y=276580 $D=21
M111 1 2 1 cpoly_p w=3.8e-06 l=2e-06 c=5.2038e-14 as=2.31158e-13 ad=7.488e-13 ps=1.44e-06 pd=1.11673e-06 sim_w=2.88e-06 m_per_maxw=1.31944 numb_sub_cont=3 nfing=1 $X=-333100 $Y=276580 $D=21
M112 1 2 1 cpoly_p w=3.8e-06 l=2e-06 c=5.2038e-14 as=2.31158e-13 ad=7.488e-13 ps=1.44e-06 pd=1.11673e-06 sim_w=2.88e-06 m_per_maxw=1.31944 numb_sub_cont=3 nfing=1 $X=-330580 $Y=276580 $D=21
M113 1 2 1 cpoly_p w=3.8e-06 l=2e-06 c=5.2038e-14 as=2.31158e-13 ad=7.488e-13 ps=1.44e-06 pd=1.11673e-06 sim_w=2.88e-06 m_per_maxw=1.31944 numb_sub_cont=3 nfing=1 $X=-328060 $Y=276580 $D=21
M114 1 2 1 cpoly_p w=3.8e-06 l=2e-06 c=5.2038e-14 as=2.31158e-13 ad=7.488e-13 ps=1.44e-06 pd=1.11673e-06 sim_w=2.88e-06 m_per_maxw=1.31944 numb_sub_cont=3 nfing=1 $X=-325540 $Y=276580 $D=21
M115 1 2 1 cpoly_p w=3.8e-06 l=2e-06 c=5.2038e-14 as=2.31158e-13 ad=7.488e-13 ps=1.44e-06 pd=1.11673e-06 sim_w=2.88e-06 m_per_maxw=1.31944 numb_sub_cont=3 nfing=1 $X=-323020 $Y=276580 $D=21
M116 1 2 1 cpoly_p w=3.8e-06 l=2e-06 c=5.2038e-14 as=2.31158e-13 ad=7.488e-13 ps=1.44e-06 pd=1.11673e-06 sim_w=2.88e-06 m_per_maxw=1.31944 numb_sub_cont=3 nfing=1 $X=-320500 $Y=276580 $D=21
M117 1 2 1 cpoly_p w=3.8e-06 l=2e-06 c=5.2038e-14 as=2.31158e-13 ad=7.488e-13 ps=1.44e-06 pd=1.11673e-06 sim_w=2.88e-06 m_per_maxw=1.31944 numb_sub_cont=3 nfing=1 $X=-317980 $Y=276580 $D=21
M118 1 2 1 cpoly_p w=3.8e-06 l=2e-06 c=5.2038e-14 as=2.31158e-13 ad=7.488e-13 ps=1.44e-06 pd=1.11673e-06 sim_w=2.88e-06 m_per_maxw=1.31944 numb_sub_cont=3 nfing=1 $X=-315460 $Y=276580 $D=21
M119 1 2 1 cpoly_p w=3.8e-06 l=2e-06 c=5.2038e-14 as=2.31158e-13 ad=7.488e-13 ps=1.44e-06 pd=1.11673e-06 sim_w=2.88e-06 m_per_maxw=1.31944 numb_sub_cont=3 nfing=1 $X=-312940 $Y=276580 $D=21
M120 1 2 1 cpoly_p w=3.8e-06 l=2e-06 c=5.2038e-14 as=2.31158e-13 ad=7.488e-13 ps=1.44e-06 pd=1.11673e-06 sim_w=2.88e-06 m_per_maxw=1.31944 numb_sub_cont=3 nfing=1 $X=-310420 $Y=276580 $D=21
M121 1 2 1 cpoly_p w=3.8e-06 l=2e-06 c=5.2038e-14 as=2.31158e-13 ad=7.488e-13 ps=1.44e-06 pd=1.11673e-06 sim_w=2.88e-06 m_per_maxw=1.31944 numb_sub_cont=3 nfing=1 $X=-307900 $Y=276580 $D=21
M122 1 2 1 cpoly_p w=3.8e-06 l=2e-06 c=5.2038e-14 as=2.31158e-13 ad=7.488e-13 ps=1.44e-06 pd=1.11673e-06 sim_w=2.88e-06 m_per_maxw=1.31944 numb_sub_cont=3 nfing=1 $X=-305380 $Y=276580 $D=21
M123 1 2 1 cpoly_p w=3.8e-06 l=2e-06 c=5.2038e-14 as=2.31158e-13 ad=7.488e-13 ps=1.44e-06 pd=1.11673e-06 sim_w=2.88e-06 m_per_maxw=1.31944 numb_sub_cont=3 nfing=1 $X=-302860 $Y=276580 $D=21
M124 1 2 1 cpoly_p w=3.8e-06 l=2e-06 c=5.2038e-14 as=2.31158e-13 ad=7.488e-13 ps=1.44e-06 pd=1.11673e-06 sim_w=2.88e-06 m_per_maxw=1.31944 numb_sub_cont=3 nfing=1 $X=-300340 $Y=276580 $D=21
M125 1 2 1 cpoly_p w=3.8e-06 l=2e-06 c=5.2038e-14 as=2.31158e-13 ad=7.488e-13 ps=1.44e-06 pd=1.11673e-06 sim_w=2.88e-06 m_per_maxw=1.31944 numb_sub_cont=3 nfing=1 $X=-297820 $Y=276580 $D=21
M126 1 2 1 cpoly_p w=3.8e-06 l=2e-06 c=5.2038e-14 as=2.31158e-13 ad=7.488e-13 ps=1.44e-06 pd=1.11673e-06 sim_w=2.88e-06 m_per_maxw=1.31944 numb_sub_cont=3 nfing=1 $X=-295300 $Y=276580 $D=21
M127 1 2 1 cpoly_p w=3.8e-06 l=2e-06 c=5.2038e-14 as=2.31158e-13 ad=7.488e-13 ps=1.44e-06 pd=1.11673e-06 sim_w=2.88e-06 m_per_maxw=1.31944 numb_sub_cont=3 nfing=1 $X=-292780 $Y=276580 $D=21
M128 1 2 1 cpoly_p w=3.8e-06 l=2e-06 c=5.2038e-14 as=2.31158e-13 ad=7.488e-13 ps=1.44e-06 pd=1.11673e-06 sim_w=2.88e-06 m_per_maxw=1.31944 numb_sub_cont=3 nfing=1 $X=-290260 $Y=276580 $D=21
M129 1 2 1 cpoly_p w=3.8e-06 l=2e-06 c=5.2038e-14 as=2.31158e-13 ad=7.488e-13 ps=1.44e-06 pd=1.11673e-06 sim_w=2.88e-06 m_per_maxw=1.31944 numb_sub_cont=3 nfing=1 $X=-287740 $Y=276580 $D=21
M130 1 2 1 cpoly_p w=3.8e-06 l=2e-06 c=5.2038e-14 as=2.31158e-13 ad=7.488e-13 ps=1.44e-06 pd=1.11673e-06 sim_w=2.88e-06 m_per_maxw=1.31944 numb_sub_cont=3 nfing=1 $X=-285220 $Y=276580 $D=21
M131 1 2 1 cpoly_p w=3.8e-06 l=2e-06 c=5.2038e-14 as=2.31158e-13 ad=7.488e-13 ps=1.44e-06 pd=1.11673e-06 sim_w=2.88e-06 m_per_maxw=1.31944 numb_sub_cont=3 nfing=1 $X=-282700 $Y=276580 $D=21
M132 1 2 1 cpoly_p w=3.8e-06 l=2e-06 c=5.2038e-14 as=2.31158e-13 ad=7.488e-13 ps=1.44e-06 pd=1.11673e-06 sim_w=2.88e-06 m_per_maxw=1.31944 numb_sub_cont=3 nfing=1 $X=-280180 $Y=276580 $D=21
M133 1 2 1 cpoly_p w=3.8e-06 l=2e-06 c=5.2038e-14 as=2.31158e-13 ad=7.488e-13 ps=1.44e-06 pd=1.11673e-06 sim_w=2.88e-06 m_per_maxw=1.31944 numb_sub_cont=3 nfing=1 $X=-277660 $Y=276580 $D=21
M134 1 2 1 cpoly_p w=3.8e-06 l=2e-06 c=5.2038e-14 as=2.31158e-13 ad=7.488e-13 ps=1.44e-06 pd=1.11673e-06 sim_w=2.88e-06 m_per_maxw=1.31944 numb_sub_cont=3 nfing=1 $X=-275140 $Y=276580 $D=21
M135 1 2 1 cpoly_p w=3.8e-06 l=2e-06 c=5.2038e-14 as=2.31158e-13 ad=7.488e-13 ps=1.44e-06 pd=1.11673e-06 sim_w=2.88e-06 m_per_maxw=1.31944 numb_sub_cont=3 nfing=1 $X=-272620 $Y=276580 $D=21
M136 1 2 1 cpoly_p w=3.8e-06 l=2e-06 c=5.2038e-14 as=2.31158e-13 ad=7.488e-13 ps=1.44e-06 pd=1.11673e-06 sim_w=2.88e-06 m_per_maxw=1.31944 numb_sub_cont=3 nfing=1 $X=-270100 $Y=276580 $D=21
M137 1 2 1 cpoly_p w=3.8e-06 l=2e-06 c=5.2038e-14 as=2.31158e-13 ad=7.488e-13 ps=1.44e-06 pd=1.11673e-06 sim_w=2.88e-06 m_per_maxw=1.31944 numb_sub_cont=3 nfing=1 $X=-267580 $Y=276580 $D=21
M138 1 2 1 cpoly_p w=3.8e-06 l=2e-06 c=5.2038e-14 as=2.31158e-13 ad=7.488e-13 ps=1.44e-06 pd=1.11673e-06 sim_w=2.88e-06 m_per_maxw=1.31944 numb_sub_cont=3 nfing=1 $X=-265060 $Y=276580 $D=21
M139 1 2 1 cpoly_p w=3.8e-06 l=2e-06 c=5.2038e-14 as=2.31158e-13 ad=7.488e-13 ps=1.44e-06 pd=1.11673e-06 sim_w=2.88e-06 m_per_maxw=1.31944 numb_sub_cont=3 nfing=1 $X=-262540 $Y=276580 $D=21
M140 1 2 1 cpoly_p w=3.8e-06 l=2e-06 c=5.2038e-14 as=2.31158e-13 ad=7.488e-13 ps=1.44e-06 pd=1.11673e-06 sim_w=2.88e-06 m_per_maxw=1.31944 numb_sub_cont=3 nfing=1 $X=-260020 $Y=276580 $D=21
M141 1 2 1 cpoly_p w=3.8e-06 l=2e-06 c=5.2038e-14 as=2.31158e-13 ad=7.488e-13 ps=1.44e-06 pd=1.11673e-06 sim_w=2.88e-06 m_per_maxw=1.31944 numb_sub_cont=3 nfing=1 $X=-257500 $Y=276580 $D=21
M142 1 2 1 cpoly_p w=3.8e-06 l=2e-06 c=5.2038e-14 as=2.31158e-13 ad=7.488e-13 ps=1.44e-06 pd=1.11673e-06 sim_w=2.88e-06 m_per_maxw=1.31944 numb_sub_cont=3 nfing=1 $X=-254980 $Y=276580 $D=21
M143 1 2 1 cpoly_p w=3.8e-06 l=2e-06 c=5.2038e-14 as=2.31158e-13 ad=7.488e-13 ps=1.44e-06 pd=1.11673e-06 sim_w=2.88e-06 m_per_maxw=1.31944 numb_sub_cont=3 nfing=1 $X=-252460 $Y=276580 $D=21
M144 1 2 1 cpoly_p w=3.8e-06 l=2e-06 c=5.2038e-14 as=2.31158e-13 ad=7.488e-13 ps=1.44e-06 pd=1.11673e-06 sim_w=2.88e-06 m_per_maxw=1.31944 numb_sub_cont=3 nfing=1 $X=-249940 $Y=276580 $D=21
M145 1 2 1 cpoly_p w=3.8e-06 l=2e-06 c=5.2038e-14 as=2.31158e-13 ad=7.488e-13 ps=1.44e-06 pd=1.11673e-06 sim_w=2.88e-06 m_per_maxw=1.31944 numb_sub_cont=3 nfing=1 $X=-247420 $Y=276580 $D=21
M146 1 2 1 cpoly_p w=3.8e-06 l=2e-06 c=5.2038e-14 as=2.31158e-13 ad=7.488e-13 ps=1.44e-06 pd=1.11673e-06 sim_w=2.88e-06 m_per_maxw=1.31944 numb_sub_cont=3 nfing=1 $X=-244900 $Y=276580 $D=21
M147 1 2 1 cpoly_p w=3.8e-06 l=2e-06 c=5.2038e-14 as=2.31158e-13 ad=7.488e-13 ps=1.44e-06 pd=1.11673e-06 sim_w=2.88e-06 m_per_maxw=1.31944 numb_sub_cont=3 nfing=1 $X=-242380 $Y=276580 $D=21
M148 1 2 1 cpoly_p w=3.8e-06 l=2e-06 c=5.2038e-14 as=2.31158e-13 ad=7.488e-13 ps=1.44e-06 pd=1.11673e-06 sim_w=2.88e-06 m_per_maxw=1.31944 numb_sub_cont=3 nfing=1 $X=-239860 $Y=276580 $D=21
M149 1 2 1 cpoly_p w=3.8e-06 l=2e-06 c=5.2038e-14 as=2.31158e-13 ad=7.488e-13 ps=1.44e-06 pd=1.11673e-06 sim_w=2.88e-06 m_per_maxw=1.31944 numb_sub_cont=3 nfing=1 $X=-237340 $Y=276580 $D=21
M150 1 2 1 cpoly_p w=3.8e-06 l=2e-06 c=5.2038e-14 as=2.31158e-13 ad=7.488e-13 ps=1.44e-06 pd=1.11673e-06 sim_w=2.88e-06 m_per_maxw=1.31944 numb_sub_cont=3 nfing=1 $X=-234820 $Y=276580 $D=21
M151 1 2 1 cpoly_p w=3.8e-06 l=2e-06 c=5.2038e-14 as=2.31158e-13 ad=7.488e-13 ps=1.44e-06 pd=1.11673e-06 sim_w=2.88e-06 m_per_maxw=1.31944 numb_sub_cont=3 nfing=1 $X=-232300 $Y=276580 $D=21
M152 1 2 1 cpoly_p w=3.8e-06 l=2e-06 c=5.2038e-14 as=2.31158e-13 ad=7.488e-13 ps=1.44e-06 pd=1.11673e-06 sim_w=2.88e-06 m_per_maxw=1.31944 numb_sub_cont=3 nfing=1 $X=-229780 $Y=276580 $D=21
M153 1 2 1 cpoly_p w=3.8e-06 l=2e-06 c=5.2038e-14 as=2.31158e-13 ad=7.488e-13 ps=1.44e-06 pd=1.11673e-06 sim_w=2.88e-06 m_per_maxw=1.31944 numb_sub_cont=3 nfing=1 $X=-227260 $Y=276580 $D=21
M154 1 2 1 cpoly_p w=3.8e-06 l=2e-06 c=5.2038e-14 as=2.31158e-13 ad=7.488e-13 ps=1.44e-06 pd=1.11673e-06 sim_w=2.88e-06 m_per_maxw=1.31944 numb_sub_cont=3 nfing=1 $X=-224740 $Y=276580 $D=21
M155 1 2 1 cpoly_p w=3.8e-06 l=2e-06 c=5.2038e-14 as=2.31158e-13 ad=7.488e-13 ps=1.44e-06 pd=1.11673e-06 sim_w=2.88e-06 m_per_maxw=1.31944 numb_sub_cont=3 nfing=1 $X=-222220 $Y=276580 $D=21
M156 1 2 1 cpoly_p w=3.8e-06 l=2e-06 c=5.2038e-14 as=2.31158e-13 ad=7.488e-13 ps=1.44e-06 pd=1.11673e-06 sim_w=2.88e-06 m_per_maxw=1.31944 numb_sub_cont=3 nfing=1 $X=-219700 $Y=276580 $D=21
M157 1 2 1 cpoly_p w=3.8e-06 l=2e-06 c=5.2038e-14 as=2.31158e-13 ad=1.152e-12 ps=1.44e-06 pd=2.23347e-06 sim_w=2.88e-06 m_per_maxw=1.31944 numb_sub_cont=3 nfing=1 $X=-217180 $Y=276580 $D=21
M158 2 1 2 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=-395880 $Y=283540 $D=22
M159 2 1 2 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=-393360 $Y=283540 $D=22
M160 2 1 2 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=-390840 $Y=283540 $D=22
M161 2 1 2 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=-388320 $Y=283540 $D=22
M162 2 1 2 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=-385800 $Y=283540 $D=22
M163 2 1 2 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=-383280 $Y=283540 $D=22
M164 2 1 2 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=-380760 $Y=283540 $D=22
M165 2 1 2 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=-378240 $Y=283540 $D=22
M166 2 1 2 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=-375720 $Y=283540 $D=22
M167 2 1 2 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=-373200 $Y=283540 $D=22
M168 2 1 2 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=-370680 $Y=283540 $D=22
M169 2 1 2 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=-368160 $Y=283540 $D=22
M170 2 1 2 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=-365640 $Y=283540 $D=22
M171 2 1 2 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=-363120 $Y=283540 $D=22
M172 2 1 2 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=-360600 $Y=283540 $D=22
M173 2 1 2 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=-358080 $Y=283540 $D=22
M174 2 1 2 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=-355560 $Y=283540 $D=22
M175 2 1 2 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=-353040 $Y=283540 $D=22
M176 2 1 2 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=-350520 $Y=283540 $D=22
M177 2 1 2 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=-348000 $Y=283540 $D=22
M178 2 1 2 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=-345480 $Y=283540 $D=22
M179 2 1 2 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=-342960 $Y=283540 $D=22
M180 2 1 2 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=-340440 $Y=283540 $D=22
M181 2 1 2 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=-337920 $Y=283540 $D=22
M182 2 1 2 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=-335400 $Y=283540 $D=22
M183 2 1 2 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=-332880 $Y=283540 $D=22
M184 2 1 2 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=-330360 $Y=283540 $D=22
M185 2 1 2 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=-327840 $Y=283540 $D=22
M186 2 1 2 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=-325320 $Y=283540 $D=22
M187 2 1 2 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=-322800 $Y=283540 $D=22
M188 2 1 2 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=-320280 $Y=283540 $D=22
M189 2 1 2 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=-317760 $Y=283540 $D=22
M190 2 1 2 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=-315240 $Y=283540 $D=22
M191 2 1 2 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=-312720 $Y=283540 $D=22
M192 2 1 2 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=-310200 $Y=283540 $D=22
M193 2 1 2 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=-307680 $Y=283540 $D=22
M194 2 1 2 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=-305160 $Y=283540 $D=22
M195 2 1 2 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=-302640 $Y=283540 $D=22
M196 2 1 2 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=-300120 $Y=283540 $D=22
M197 2 1 2 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=-297600 $Y=283540 $D=22
M198 2 1 2 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=-295080 $Y=283540 $D=22
M199 2 1 2 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=-292560 $Y=283540 $D=22
M200 2 1 2 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=-290040 $Y=283540 $D=22
M201 2 1 2 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=-287520 $Y=283540 $D=22
M202 2 1 2 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=-285000 $Y=283540 $D=22
M203 2 1 2 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=-282480 $Y=283540 $D=22
M204 2 1 2 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=-279960 $Y=283540 $D=22
M205 2 1 2 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=-277440 $Y=283540 $D=22
M206 2 1 2 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=-274920 $Y=283540 $D=22
M207 2 1 2 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=-272400 $Y=283540 $D=22
M208 2 1 2 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=-269880 $Y=283540 $D=22
M209 2 1 2 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=-267360 $Y=283540 $D=22
M210 2 1 2 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=-264840 $Y=283540 $D=22
M211 2 1 2 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=-262320 $Y=283540 $D=22
M212 2 1 2 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=-259800 $Y=283540 $D=22
M213 2 1 2 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=-257280 $Y=283540 $D=22
M214 2 1 2 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=-254760 $Y=283540 $D=22
M215 2 1 2 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=-252240 $Y=283540 $D=22
M216 2 1 2 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=-249720 $Y=283540 $D=22
M217 2 1 2 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=-247200 $Y=283540 $D=22
M218 2 1 2 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=-244680 $Y=283540 $D=22
M219 2 1 2 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=-242160 $Y=283540 $D=22
M220 2 1 2 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=-239640 $Y=283540 $D=22
M221 2 1 2 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=-237120 $Y=283540 $D=22
M222 2 1 2 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=-234600 $Y=283540 $D=22
M223 2 1 2 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=-232080 $Y=283540 $D=22
M224 2 1 2 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=-229560 $Y=283540 $D=22
M225 2 1 2 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=-227040 $Y=283540 $D=22
M226 2 1 2 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=-224520 $Y=283540 $D=22
M227 2 1 2 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=-222000 $Y=283540 $D=22
M228 2 1 2 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=-219480 $Y=283540 $D=22
M229 2 1 2 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=-216960 $Y=283540 $D=22
M230 2 1 2 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=-214440 $Y=283540 $D=22
M231 2 1 2 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=-211920 $Y=283540 $D=22
M232 2 1 2 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=-209400 $Y=283540 $D=22
M233 2 1 2 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=-206880 $Y=283540 $D=22
M234 2 1 2 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=-204360 $Y=283540 $D=22
M235 2 1 2 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=-201840 $Y=283540 $D=22
M236 2 1 2 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=-199320 $Y=283540 $D=22
X293 7 8 17 18 ICV_150 $T=-395840 271760 1 0 $X=-396200 $Y=268540
X294 7 8 17 18 ICV_150 $T=-395840 271760 0 0 $X=-396200 $Y=271420
X295 7 8 17 18 ICV_150 $T=-371680 271760 1 0 $X=-372040 $Y=268540
X296 7 8 17 18 ICV_150 $T=-371680 271760 0 0 $X=-372040 $Y=271420
X297 7 8 17 18 ICV_150 $T=-347520 271760 1 0 $X=-347880 $Y=268540
X298 7 8 17 18 ICV_150 $T=-347520 271760 0 0 $X=-347880 $Y=271420
X299 7 8 17 18 ICV_150 $T=-323360 271760 1 0 $X=-323720 $Y=268540
X300 7 8 17 18 ICV_150 $T=-323360 271760 0 0 $X=-323720 $Y=271420
X301 7 8 17 18 ICV_150 $T=-299200 271760 1 0 $X=-299560 $Y=268540
X302 7 8 17 18 ICV_150 $T=-299200 271760 0 0 $X=-299560 $Y=271420
X303 7 8 17 18 ICV_150 $T=-275040 271760 1 0 $X=-275400 $Y=268540
X304 7 8 17 18 ICV_150 $T=-275040 271760 0 0 $X=-275400 $Y=271420
X305 7 8 17 18 ICV_150 $T=-250880 271760 1 0 $X=-251240 $Y=268540
X306 7 8 17 18 ICV_150 $T=-250880 271760 0 0 $X=-251240 $Y=271420
.ENDS
***************************************
.SUBCKT pmos_a_CDNS_5887047866539 1 2 3
** N=3 EP=3 IP=0 FDC=1
M0 2 3 1 1 pmos_a L=3e-07 W=1.2e-06 AD=7.2e-13 AS=1.62e-13 PD=1.8e-06 PS=9e-07 w_cont=6e-07 nfing=1 mmm=1 $X=620 $Y=200 $D=5
.ENDS
***************************************
.SUBCKT ICV_152 1 2 3 4 5 6 7 9 10 11 12 15
** N=16 EP=12 IP=140 FDC=88
*.SEEDPROM
M0 5 15 5 5 nmos_a L=2e-06 W=9.26e-05 AD=7.90041e-13 AS=2.4076e-11 PD=1.51931e-06 PS=1.51931e-06 w_cont=5.1e-06 nfing=1 source_num=2 $X=-200600 $Y=160080 $D=1
M1 5 15 5 5 nmos_a L=2e-06 W=9.26e-05 AD=7.90041e-13 AS=3.704e-11 PD=1.51931e-06 PS=1.51931e-06 w_cont=5.1e-06 nfing=1 source_num=2 $X=-198080 $Y=160080 $D=1
M2 5 15 5 5 nmos_a L=2e-06 W=9.26e-05 AD=7.90041e-13 AS=3.704e-11 PD=1.51931e-06 PS=1.51931e-06 w_cont=5.1e-06 nfing=1 source_num=2 $X=-311480 $Y=160080 $D=1
M3 5 15 5 5 nmos_a L=2e-06 W=9.26e-05 AD=7.90041e-13 AS=2.4076e-11 PD=1.51931e-06 PS=1.51931e-06 w_cont=5.1e-06 nfing=1 source_num=2 $X=-301400 $Y=160080 $D=1
M4 5 15 5 5 nmos_a L=2e-06 W=9.26e-05 AD=7.90041e-13 AS=2.4076e-11 PD=1.51931e-06 PS=1.51931e-06 w_cont=5.1e-06 nfing=1 source_num=2 $X=-291320 $Y=160080 $D=1
M5 5 15 5 5 nmos_a L=2e-06 W=9.26e-05 AD=7.90041e-13 AS=2.4076e-11 PD=1.51931e-06 PS=1.51931e-06 w_cont=5.1e-06 nfing=1 source_num=2 $X=-281240 $Y=160080 $D=1
M6 5 15 5 5 nmos_a L=2e-06 W=9.26e-05 AD=7.90041e-13 AS=2.4076e-11 PD=1.51931e-06 PS=1.51931e-06 w_cont=5.1e-06 nfing=1 source_num=2 $X=-271160 $Y=160080 $D=1
M7 5 15 5 5 nmos_a L=2e-06 W=9.26e-05 AD=7.90041e-13 AS=2.4076e-11 PD=1.51931e-06 PS=1.51931e-06 w_cont=5.1e-06 nfing=1 source_num=2 $X=-261080 $Y=160080 $D=1
M8 5 15 5 5 nmos_a L=2e-06 W=9.26e-05 AD=7.90041e-13 AS=2.4076e-11 PD=1.51931e-06 PS=1.51931e-06 w_cont=5.1e-06 nfing=1 source_num=2 $X=-251000 $Y=160080 $D=1
M9 5 15 5 5 nmos_a L=2e-06 W=9.26e-05 AD=7.90041e-13 AS=2.4076e-11 PD=1.51931e-06 PS=1.51931e-06 w_cont=5.1e-06 nfing=1 source_num=2 $X=-240920 $Y=160080 $D=1
M10 5 15 5 5 nmos_a L=2e-06 W=9.26e-05 AD=7.90041e-13 AS=2.4076e-11 PD=1.51931e-06 PS=1.51931e-06 w_cont=5.1e-06 nfing=1 source_num=2 $X=-230840 $Y=160080 $D=1
M11 5 15 5 5 nmos_a L=2e-06 W=9.26e-05 AD=7.90041e-13 AS=2.4076e-11 PD=1.51931e-06 PS=1.51931e-06 w_cont=5.1e-06 nfing=1 source_num=2 $X=-220760 $Y=160080 $D=1
M12 5 15 5 5 nmos_a L=2e-06 W=9.26e-05 AD=7.90041e-13 AS=2.4076e-11 PD=1.51931e-06 PS=1.51931e-06 w_cont=5.1e-06 nfing=1 source_num=2 $X=-210680 $Y=160080 $D=1
M13 6 7 1 1 nmos_a L=3e-07 W=4.8e-07 AD=2.808e-13 AS=1.92e-13 PD=5.4e-07 PS=5.4e-07 w_cont=6e-07 nfing=1 source_num=2 $X=-223460 $Y=265260 $D=1
M14 6 7 1 1 nmos_a L=3e-07 W=4.8e-07 AD=2.808e-13 AS=1.92e-13 PD=5.4e-07 PS=5.4e-07 w_cont=6e-07 nfing=1 source_num=2 $X=-223460 $Y=266740 $D=1
M15 6 7 1 1 nmos_a L=3e-07 W=4.8e-07 AD=2.808e-13 AS=1.248e-13 PD=5.4e-07 PS=5.4e-07 w_cont=6e-07 nfing=1 source_num=2 $X=-222640 $Y=265260 $D=1
M16 6 7 1 1 nmos_a L=3e-07 W=4.8e-07 AD=2.808e-13 AS=1.248e-13 PD=5.4e-07 PS=5.4e-07 w_cont=6e-07 nfing=1 source_num=2 $X=-222640 $Y=266740 $D=1
M17 7 7 1 1 nmos_a L=3e-07 W=4.8e-07 AD=2.808e-13 AS=1.248e-13 PD=5.4e-07 PS=5.4e-07 w_cont=6e-07 nfing=1 source_num=2 $X=-221820 $Y=265260 $D=1
M18 6 7 1 1 nmos_a L=3e-07 W=4.8e-07 AD=2.808e-13 AS=1.248e-13 PD=5.4e-07 PS=5.4e-07 w_cont=6e-07 nfing=1 source_num=2 $X=-221820 $Y=266740 $D=1
M19 7 7 1 1 nmos_a L=3e-07 W=4.8e-07 AD=2.808e-13 AS=1.248e-13 PD=5.4e-07 PS=5.4e-07 w_cont=6e-07 nfing=1 source_num=2 $X=-221000 $Y=265260 $D=1
M20 6 7 1 1 nmos_a L=3e-07 W=4.8e-07 AD=2.808e-13 AS=1.248e-13 PD=5.4e-07 PS=5.4e-07 w_cont=6e-07 nfing=1 source_num=2 $X=-221000 $Y=266740 $D=1
M21 6 7 1 1 nmos_a L=3e-07 W=4.8e-07 AD=2.808e-13 AS=1.248e-13 PD=5.4e-07 PS=5.4e-07 w_cont=6e-07 nfing=1 source_num=2 $X=-220180 $Y=265260 $D=1
M22 6 7 1 1 nmos_a L=3e-07 W=4.8e-07 AD=2.808e-13 AS=1.248e-13 PD=5.4e-07 PS=5.4e-07 w_cont=6e-07 nfing=1 source_num=2 $X=-220180 $Y=266740 $D=1
M23 6 7 1 1 nmos_a L=3e-07 W=4.8e-07 AD=2.808e-13 AS=1.248e-13 PD=5.4e-07 PS=5.4e-07 w_cont=6e-07 nfing=1 source_num=2 $X=-219360 $Y=265260 $D=1
M24 6 7 1 1 nmos_a L=3e-07 W=4.8e-07 AD=2.808e-13 AS=1.248e-13 PD=5.4e-07 PS=5.4e-07 w_cont=6e-07 nfing=1 source_num=2 $X=-219360 $Y=266740 $D=1
M25 7 7 1 1 nmos_a L=3e-07 W=4.8e-07 AD=2.808e-13 AS=1.248e-13 PD=5.4e-07 PS=5.4e-07 w_cont=6e-07 nfing=1 source_num=2 $X=-218540 $Y=265260 $D=1
M26 6 7 1 1 nmos_a L=3e-07 W=4.8e-07 AD=2.808e-13 AS=1.248e-13 PD=5.4e-07 PS=5.4e-07 w_cont=6e-07 nfing=1 source_num=2 $X=-218540 $Y=266740 $D=1
M27 7 7 1 1 nmos_a L=3e-07 W=4.8e-07 AD=2.808e-13 AS=1.248e-13 PD=5.4e-07 PS=5.4e-07 w_cont=6e-07 nfing=1 source_num=2 $X=-217720 $Y=265260 $D=1
M28 6 7 1 1 nmos_a L=3e-07 W=4.8e-07 AD=2.808e-13 AS=1.248e-13 PD=5.4e-07 PS=5.4e-07 w_cont=6e-07 nfing=1 source_num=2 $X=-217720 $Y=266740 $D=1
M29 6 7 1 1 nmos_a L=3e-07 W=4.8e-07 AD=2.808e-13 AS=1.248e-13 PD=5.4e-07 PS=5.4e-07 w_cont=6e-07 nfing=1 source_num=2 $X=-216900 $Y=265260 $D=1
M30 6 7 1 1 nmos_a L=3e-07 W=4.8e-07 AD=2.808e-13 AS=1.248e-13 PD=5.4e-07 PS=5.4e-07 w_cont=6e-07 nfing=1 source_num=2 $X=-216900 $Y=266740 $D=1
M31 6 7 1 1 nmos_a L=3e-07 W=4.8e-07 AD=2.808e-13 AS=1.92e-13 PD=5.4e-07 PS=5.4e-07 w_cont=6e-07 nfing=1 source_num=2 $X=-216080 $Y=265260 $D=1
M32 6 7 1 1 nmos_a L=3e-07 W=4.8e-07 AD=2.808e-13 AS=1.92e-13 PD=5.4e-07 PS=5.4e-07 w_cont=6e-07 nfing=1 source_num=2 $X=-216080 $Y=266740 $D=1
M33 11 10 2 2 pmos_a L=2.4e-07 W=4.8e-07 AD=4.32e-13 AS=1.224e-13 PD=1.08e-06 PS=5.4e-07 w_cont=6e-07 nfing=1 mmm=1 $X=-200580 $Y=267560 $D=5
M34 12 10 2 2 pmos_a L=2.4e-07 W=4.8e-07 AD=4.32e-13 AS=1.224e-13 PD=1.08e-06 PS=5.4e-07 w_cont=6e-07 nfing=1 mmm=1 $X=-199100 $Y=267560 $D=5
R35 2 3 108140 L=0.0001605 W=5e-07 m=1 $[rppoly] $X=-385280 $Y=261340 $D=19
X36 1 5 10 nmos_a_CDNS_5887047866553 $T=-293080 259920 0 270 $X=-293080 $Y=258480
X37 1 5 10 nmos_a_CDNS_5887047866553 $T=-273680 259920 0 270 $X=-273680 $Y=258480
X38 1 5 10 nmos_a_CDNS_5887047866553 $T=-254120 259920 0 270 $X=-254120 $Y=258480
X39 1 5 10 nmos_a_CDNS_5887047866553 $T=-234720 259920 0 270 $X=-234720 $Y=258480
X40 1 5 10 nmos_a_CDNS_5887047866553 $T=-214940 259920 0 270 $X=-214940 $Y=258480
X42 5 15 ICV_135 $T=-312100 159880 0 0 $X=-312100 $Y=159880
X43 5 15 ICV_135 $T=-302020 159880 0 0 $X=-302020 $Y=159880
X44 5 15 ICV_135 $T=-291940 159880 0 0 $X=-291940 $Y=159880
X45 5 15 ICV_135 $T=-281860 159880 0 0 $X=-281860 $Y=159880
X46 5 15 ICV_135 $T=-271780 159880 0 0 $X=-271780 $Y=159880
X47 5 15 ICV_135 $T=-261700 159880 0 0 $X=-261700 $Y=159880
X48 5 15 ICV_135 $T=-251620 159880 0 0 $X=-251620 $Y=159880
X49 5 15 ICV_135 $T=-241540 159880 0 0 $X=-241540 $Y=159880
X50 5 15 ICV_135 $T=-231460 159880 0 0 $X=-231460 $Y=159880
X51 5 15 ICV_135 $T=-221380 159880 0 0 $X=-221380 $Y=159880
X52 5 15 ICV_135 $T=-211300 159880 0 0 $X=-211300 $Y=159880
X53 2 5 10 pmos_a_CDNS_5887047866552 $T=-293580 258480 0 90 $X=-304680 $Y=258480
X54 2 5 10 pmos_a_CDNS_5887047866552 $T=-274180 258480 0 90 $X=-285280 $Y=258480
X55 2 5 10 pmos_a_CDNS_5887047866552 $T=-254780 258480 0 90 $X=-265880 $Y=258480
X56 2 5 10 pmos_a_CDNS_5887047866552 $T=-235220 258480 0 90 $X=-246320 $Y=258480
X57 2 5 10 pmos_a_CDNS_5887047866552 $T=-215700 258480 0 90 $X=-226800 $Y=258480
X58 2 11 pmos_a_CDNS_5887047866541 $T=-203000 264940 0 0 $X=-203000 $Y=264940
X79 2 9 9 pmos_a_CDNS_5887047866539 $T=-212100 265360 1 180 $X=-213600 $Y=265360
X80 2 4 9 pmos_a_CDNS_5887047866539 $T=-212820 265360 0 0 $X=-212820 $Y=265360
X81 2 9 9 pmos_a_CDNS_5887047866539 $T=-209780 265360 1 180 $X=-211280 $Y=265360
X82 2 4 9 pmos_a_CDNS_5887047866539 $T=-210500 265360 0 0 $X=-210500 $Y=265360
X83 2 9 9 pmos_a_CDNS_5887047866539 $T=-207460 265360 1 180 $X=-208960 $Y=265360
X84 2 4 9 pmos_a_CDNS_5887047866539 $T=-208180 265360 0 0 $X=-208180 $Y=265360
X85 2 9 9 pmos_a_CDNS_5887047866539 $T=-205140 265360 1 180 $X=-206640 $Y=265360
X86 2 4 9 pmos_a_CDNS_5887047866539 $T=-205860 265360 0 0 $X=-205860 $Y=265360
.ENDS
***************************************
.SUBCKT ICV_153 3 4
** N=4 EP=2 IP=24 FDC=46
*.SEEDPROM
M0 3 4 3 3 nmos_a L=2e-06 W=9.26e-05 AD=1.21545e-12 AS=2.4076e-11 PD=3.03862e-06 PS=1.51931e-06 w_cont=5.1e-06 nfing=1 source_num=2 $X=-198080 $Y=61480 $D=1
M1 3 4 3 3 nmos_a L=2e-06 W=9.26e-05 AD=7.90041e-13 AS=2.4076e-11 PD=1.51931e-06 PS=1.51931e-06 w_cont=5.1e-06 nfing=1 source_num=2 $X=-200600 $Y=61480 $D=1
M2 3 4 3 3 nmos_a L=2e-06 W=9.26e-05 AD=1.21545e-12 AS=2.4076e-11 PD=3.03862e-06 PS=1.51931e-06 w_cont=5.1e-06 nfing=1 source_num=2 $X=-311480 $Y=61480 $D=1
M3 3 4 3 3 nmos_a L=2e-06 W=9.26e-05 AD=7.90041e-13 AS=2.4076e-11 PD=1.51931e-06 PS=1.51931e-06 w_cont=5.1e-06 nfing=1 source_num=2 $X=-301400 $Y=61480 $D=1
M4 3 4 3 3 nmos_a L=2e-06 W=9.26e-05 AD=7.90041e-13 AS=2.4076e-11 PD=1.51931e-06 PS=1.51931e-06 w_cont=5.1e-06 nfing=1 source_num=2 $X=-291320 $Y=61480 $D=1
M5 3 4 3 3 nmos_a L=2e-06 W=9.26e-05 AD=7.90041e-13 AS=2.4076e-11 PD=1.51931e-06 PS=1.51931e-06 w_cont=5.1e-06 nfing=1 source_num=2 $X=-281240 $Y=61480 $D=1
M6 3 4 3 3 nmos_a L=2e-06 W=9.26e-05 AD=7.90041e-13 AS=2.4076e-11 PD=1.51931e-06 PS=1.51931e-06 w_cont=5.1e-06 nfing=1 source_num=2 $X=-271160 $Y=61480 $D=1
M7 3 4 3 3 nmos_a L=2e-06 W=9.26e-05 AD=7.90041e-13 AS=2.4076e-11 PD=1.51931e-06 PS=1.51931e-06 w_cont=5.1e-06 nfing=1 source_num=2 $X=-261080 $Y=61480 $D=1
M8 3 4 3 3 nmos_a L=2e-06 W=9.26e-05 AD=7.90041e-13 AS=2.4076e-11 PD=1.51931e-06 PS=1.51931e-06 w_cont=5.1e-06 nfing=1 source_num=2 $X=-251000 $Y=61480 $D=1
M9 3 4 3 3 nmos_a L=2e-06 W=9.26e-05 AD=7.90041e-13 AS=2.4076e-11 PD=1.51931e-06 PS=1.51931e-06 w_cont=5.1e-06 nfing=1 source_num=2 $X=-240920 $Y=61480 $D=1
M10 3 4 3 3 nmos_a L=2e-06 W=9.26e-05 AD=7.90041e-13 AS=2.4076e-11 PD=1.51931e-06 PS=1.51931e-06 w_cont=5.1e-06 nfing=1 source_num=2 $X=-230840 $Y=61480 $D=1
M11 3 4 3 3 nmos_a L=2e-06 W=9.26e-05 AD=7.90041e-13 AS=2.4076e-11 PD=1.51931e-06 PS=1.51931e-06 w_cont=5.1e-06 nfing=1 source_num=2 $X=-220760 $Y=61480 $D=1
M12 3 4 3 3 nmos_a L=2e-06 W=9.26e-05 AD=7.90041e-13 AS=2.4076e-11 PD=1.51931e-06 PS=1.51931e-06 w_cont=5.1e-06 nfing=1 source_num=2 $X=-210680 $Y=61480 $D=1
X14 3 4 ICV_138 $T=-308860 61280 1 180 $X=-312060 $Y=61280
X15 3 4 ICV_138 $T=-298780 61280 1 180 $X=-301980 $Y=61280
X16 3 4 ICV_138 $T=-288700 61280 1 180 $X=-291900 $Y=61280
X17 3 4 ICV_138 $T=-278620 61280 1 180 $X=-281820 $Y=61280
X18 3 4 ICV_138 $T=-268540 61280 1 180 $X=-271740 $Y=61280
X19 3 4 ICV_138 $T=-258460 61280 1 180 $X=-261660 $Y=61280
X20 3 4 ICV_138 $T=-248380 61280 1 180 $X=-251580 $Y=61280
X21 3 4 ICV_138 $T=-238300 61280 1 180 $X=-241500 $Y=61280
X22 3 4 ICV_138 $T=-228220 61280 1 180 $X=-231420 $Y=61280
X23 3 4 ICV_138 $T=-218140 61280 1 180 $X=-221340 $Y=61280
X24 3 4 ICV_138 $T=-208060 61280 1 180 $X=-211260 $Y=61280
.ENDS
***************************************
.SUBCKT ICV_154 2 4 5 6 7 8 9 10 11 12
** N=12 EP=10 IP=72 FDC=100
*.SEEDPROM
M0 12 7 12 12 nmos_a L=2e-06 W=7e-05 AD=1.21125e-12 AS=1.82e-11 PD=3.02811e-06 PS=1.51406e-06 w_cont=3.6e-06 nfing=1 source_num=2 $X=-198080 $Y=-15340 $D=1
M1 12 7 12 12 nmos_a L=2e-06 W=7e-05 AD=7.8731e-13 AS=1.82e-11 PD=1.51406e-06 PS=1.51406e-06 w_cont=3.6e-06 nfing=1 source_num=2 $X=-200600 $Y=-15340 $D=1
M2 11 6 11 11 nmos_a L=2e-06 W=1.5e-05 AD=1.23648e-12 AS=3.9e-12 PD=3.0912e-06 PS=1.5456e-06 w_cont=1.1e-06 nfing=1 source_num=2 $X=-198080 $Y=-34660 $D=1
M3 11 6 11 11 nmos_a L=2e-06 W=1.5e-05 AD=8.03712e-13 AS=3.9e-12 PD=1.5456e-06 PS=1.5456e-06 w_cont=1.1e-06 nfing=1 source_num=2 $X=-200600 $Y=-34660 $D=1
M4 12 7 12 12 nmos_a L=2e-06 W=7e-05 AD=1.21125e-12 AS=1.82e-11 PD=3.02811e-06 PS=1.51406e-06 w_cont=3.6e-06 nfing=1 source_num=2 $X=-311480 $Y=-15340 $D=1
M5 12 7 12 12 nmos_a L=2e-06 W=7e-05 AD=7.8731e-13 AS=1.82e-11 PD=1.51406e-06 PS=1.51406e-06 w_cont=3.6e-06 nfing=1 source_num=2 $X=-301400 $Y=-15340 $D=1
M6 12 7 12 12 nmos_a L=2e-06 W=7e-05 AD=7.8731e-13 AS=1.82e-11 PD=1.51406e-06 PS=1.51406e-06 w_cont=3.6e-06 nfing=1 source_num=2 $X=-291320 $Y=-15340 $D=1
M7 12 7 12 12 nmos_a L=2e-06 W=7e-05 AD=7.8731e-13 AS=1.82e-11 PD=1.51406e-06 PS=1.51406e-06 w_cont=3.6e-06 nfing=1 source_num=2 $X=-281240 $Y=-15340 $D=1
M8 12 7 12 12 nmos_a L=2e-06 W=7e-05 AD=7.8731e-13 AS=1.82e-11 PD=1.51406e-06 PS=1.51406e-06 w_cont=3.6e-06 nfing=1 source_num=2 $X=-271160 $Y=-15340 $D=1
M9 12 7 12 12 nmos_a L=2e-06 W=7e-05 AD=7.8731e-13 AS=1.82e-11 PD=1.51406e-06 PS=1.51406e-06 w_cont=3.6e-06 nfing=1 source_num=2 $X=-261080 $Y=-15340 $D=1
M10 12 7 12 12 nmos_a L=2e-06 W=7e-05 AD=7.8731e-13 AS=1.82e-11 PD=1.51406e-06 PS=1.51406e-06 w_cont=3.6e-06 nfing=1 source_num=2 $X=-251000 $Y=-15340 $D=1
M11 12 7 12 12 nmos_a L=2e-06 W=7e-05 AD=7.8731e-13 AS=1.82e-11 PD=1.51406e-06 PS=1.51406e-06 w_cont=3.6e-06 nfing=1 source_num=2 $X=-240920 $Y=-15340 $D=1
M12 12 7 12 12 nmos_a L=2e-06 W=7e-05 AD=7.8731e-13 AS=1.82e-11 PD=1.51406e-06 PS=1.51406e-06 w_cont=3.6e-06 nfing=1 source_num=2 $X=-230840 $Y=-15340 $D=1
M13 12 7 12 12 nmos_a L=2e-06 W=7e-05 AD=7.8731e-13 AS=1.82e-11 PD=1.51406e-06 PS=1.51406e-06 w_cont=3.6e-06 nfing=1 source_num=2 $X=-220760 $Y=-15340 $D=1
M14 12 7 12 12 nmos_a L=2e-06 W=7e-05 AD=7.8731e-13 AS=1.82e-11 PD=1.51406e-06 PS=1.51406e-06 w_cont=3.6e-06 nfing=1 source_num=2 $X=-210680 $Y=-15340 $D=1
M15 11 6 11 11 nmos_a L=2e-06 W=1.5e-05 AD=1.23648e-12 AS=3.9e-12 PD=3.0912e-06 PS=1.5456e-06 w_cont=1.1e-06 nfing=1 source_num=2 $X=-311480 $Y=-34660 $D=1
M16 11 6 11 11 nmos_a L=2e-06 W=1.5e-05 AD=8.03712e-13 AS=3.9e-12 PD=1.5456e-06 PS=1.5456e-06 w_cont=1.1e-06 nfing=1 source_num=2 $X=-301400 $Y=-34660 $D=1
M17 11 6 11 11 nmos_a L=2e-06 W=1.5e-05 AD=8.03712e-13 AS=3.9e-12 PD=1.5456e-06 PS=1.5456e-06 w_cont=1.1e-06 nfing=1 source_num=2 $X=-291320 $Y=-34660 $D=1
M18 11 6 11 11 nmos_a L=2e-06 W=1.5e-05 AD=8.03712e-13 AS=3.9e-12 PD=1.5456e-06 PS=1.5456e-06 w_cont=1.1e-06 nfing=1 source_num=2 $X=-281240 $Y=-34660 $D=1
M19 11 6 11 11 nmos_a L=2e-06 W=1.5e-05 AD=8.03712e-13 AS=3.9e-12 PD=1.5456e-06 PS=1.5456e-06 w_cont=1.1e-06 nfing=1 source_num=2 $X=-271160 $Y=-34660 $D=1
M20 11 6 11 11 nmos_a L=2e-06 W=1.5e-05 AD=8.03712e-13 AS=3.9e-12 PD=1.5456e-06 PS=1.5456e-06 w_cont=1.1e-06 nfing=1 source_num=2 $X=-261080 $Y=-34660 $D=1
M21 11 6 11 11 nmos_a L=2e-06 W=1.5e-05 AD=8.03712e-13 AS=3.9e-12 PD=1.5456e-06 PS=1.5456e-06 w_cont=1.1e-06 nfing=1 source_num=2 $X=-251000 $Y=-34660 $D=1
M22 11 6 11 11 nmos_a L=2e-06 W=1.5e-05 AD=8.03712e-13 AS=3.9e-12 PD=1.5456e-06 PS=1.5456e-06 w_cont=1.1e-06 nfing=1 source_num=2 $X=-240920 $Y=-34660 $D=1
M23 11 6 11 11 nmos_a L=2e-06 W=1.5e-05 AD=8.03712e-13 AS=3.9e-12 PD=1.5456e-06 PS=1.5456e-06 w_cont=1.1e-06 nfing=1 source_num=2 $X=-230840 $Y=-34660 $D=1
M24 11 6 11 11 nmos_a L=2e-06 W=1.5e-05 AD=8.03712e-13 AS=3.9e-12 PD=1.5456e-06 PS=1.5456e-06 w_cont=1.1e-06 nfing=1 source_num=2 $X=-220760 $Y=-34660 $D=1
M25 11 6 11 11 nmos_a L=2e-06 W=1.5e-05 AD=8.03712e-13 AS=3.9e-12 PD=1.5456e-06 PS=1.5456e-06 w_cont=1.1e-06 nfing=1 source_num=2 $X=-210680 $Y=-34660 $D=1
X26 4 12 9 nmos_a_CDNS_5887047866553 $T=-222780 58960 1 90 $X=-222780 $Y=58960
X27 5 11 7 nmos_a_CDNS_5887047866553 $T=-208180 -17860 0 90 $X=-215480 $Y=-17860
X28 4 12 9 nmos_a_CDNS_5887047866553 $T=-203380 58960 1 90 $X=-203380 $Y=58960
X29 2 12 9 pmos_a_CDNS_5887047866552 $T=-223280 60440 1 270 $X=-234380 $Y=59000
X30 2 12 9 pmos_a_CDNS_5887047866552 $T=-203880 60440 1 270 $X=-214980 $Y=59000
X31 4 11 7 pmos_a_CDNS_5887047866552 $T=-207680 -16380 0 270 $X=-207680 $Y=-17820
X34 12 7 ICV_142 $T=-308860 -15540 1 180 $X=-312060 $Y=-15540
X35 12 7 ICV_142 $T=-298780 -15540 1 180 $X=-301980 $Y=-15540
X36 12 7 ICV_142 $T=-288700 -15540 1 180 $X=-291900 $Y=-15540
X37 12 7 ICV_142 $T=-278620 -15540 1 180 $X=-281820 $Y=-15540
X38 12 7 ICV_142 $T=-268540 -15540 1 180 $X=-271740 $Y=-15540
X39 12 7 ICV_142 $T=-258460 -15540 1 180 $X=-261660 $Y=-15540
X40 12 7 ICV_142 $T=-248380 -15540 1 180 $X=-251580 $Y=-15540
X41 12 7 ICV_142 $T=-238300 -15540 1 180 $X=-241500 $Y=-15540
X42 12 7 ICV_142 $T=-228220 -15540 1 180 $X=-231420 $Y=-15540
X43 12 7 ICV_142 $T=-218140 -15540 1 180 $X=-221340 $Y=-15540
X44 12 7 ICV_142 $T=-208060 -15540 1 180 $X=-211260 $Y=-15540
X45 11 6 ICV_143 $T=-308860 -34860 1 180 $X=-312060 $Y=-34860
X46 11 6 ICV_143 $T=-298780 -34860 1 180 $X=-301980 $Y=-34860
X47 11 6 ICV_143 $T=-288700 -34860 1 180 $X=-291900 $Y=-34860
X48 11 6 ICV_143 $T=-278620 -34860 1 180 $X=-281820 $Y=-34860
X49 11 6 ICV_143 $T=-268540 -34860 1 180 $X=-271740 $Y=-34860
X50 11 6 ICV_143 $T=-258460 -34860 1 180 $X=-261660 $Y=-34860
X51 11 6 ICV_143 $T=-248380 -34860 1 180 $X=-251580 $Y=-34860
X52 11 6 ICV_143 $T=-238300 -34860 1 180 $X=-241500 $Y=-34860
X53 11 6 ICV_143 $T=-228220 -34860 1 180 $X=-231420 $Y=-34860
X54 11 6 ICV_143 $T=-218140 -34860 1 180 $X=-221340 $Y=-34860
X55 11 6 ICV_143 $T=-208060 -34860 1 180 $X=-211260 $Y=-34860
X56 8 10 6 nmos_a_CDNS_5887047866558 $T=-204140 -37180 0 90 $X=-208040 $Y=-37180
X57 5 10 6 pmos_a_CDNS_5887047866557 $T=-203640 -37180 1 90 $X=-203640 $Y=-37180
.ENDS
***************************************
.SUBCKT ICV_155 4 6
** N=6 EP=2 IP=24 FDC=46
*.SEEDPROM
M0 4 6 4 4 nmos_a L=2e-06 W=0.0001 AD=1.21075e-12 AS=2.6e-11 PD=3.02688e-06 PS=1.51344e-06 w_cont=5.1e-06 nfing=1 source_num=2 $X=-198080 $Y=-142980 $D=1
M1 4 6 4 4 nmos_a L=2e-06 W=0.0001 AD=7.86989e-13 AS=2.6e-11 PD=1.51344e-06 PS=1.51344e-06 w_cont=5.1e-06 nfing=1 source_num=2 $X=-200600 $Y=-142980 $D=1
M2 4 6 4 4 nmos_a L=2e-06 W=0.0001 AD=1.21075e-12 AS=2.6e-11 PD=3.02688e-06 PS=1.51344e-06 w_cont=5.1e-06 nfing=1 source_num=2 $X=-311480 $Y=-142980 $D=1
M3 4 6 4 4 nmos_a L=2e-06 W=0.0001 AD=7.86989e-13 AS=2.6e-11 PD=1.51344e-06 PS=1.51344e-06 w_cont=5.1e-06 nfing=1 source_num=2 $X=-301400 $Y=-142980 $D=1
M4 4 6 4 4 nmos_a L=2e-06 W=0.0001 AD=7.86989e-13 AS=2.6e-11 PD=1.51344e-06 PS=1.51344e-06 w_cont=5.1e-06 nfing=1 source_num=2 $X=-291320 $Y=-142980 $D=1
M5 4 6 4 4 nmos_a L=2e-06 W=0.0001 AD=7.86989e-13 AS=2.6e-11 PD=1.51344e-06 PS=1.51344e-06 w_cont=5.1e-06 nfing=1 source_num=2 $X=-281240 $Y=-142980 $D=1
M6 4 6 4 4 nmos_a L=2e-06 W=0.0001 AD=7.86989e-13 AS=2.6e-11 PD=1.51344e-06 PS=1.51344e-06 w_cont=5.1e-06 nfing=1 source_num=2 $X=-271160 $Y=-142980 $D=1
M7 4 6 4 4 nmos_a L=2e-06 W=0.0001 AD=7.86989e-13 AS=2.6e-11 PD=1.51344e-06 PS=1.51344e-06 w_cont=5.1e-06 nfing=1 source_num=2 $X=-261080 $Y=-142980 $D=1
M8 4 6 4 4 nmos_a L=2e-06 W=0.0001 AD=7.86989e-13 AS=2.6e-11 PD=1.51344e-06 PS=1.51344e-06 w_cont=5.1e-06 nfing=1 source_num=2 $X=-251000 $Y=-142980 $D=1
M9 4 6 4 4 nmos_a L=2e-06 W=0.0001 AD=7.86989e-13 AS=2.6e-11 PD=1.51344e-06 PS=1.51344e-06 w_cont=5.1e-06 nfing=1 source_num=2 $X=-240920 $Y=-142980 $D=1
M10 4 6 4 4 nmos_a L=2e-06 W=0.0001 AD=7.86989e-13 AS=2.6e-11 PD=1.51344e-06 PS=1.51344e-06 w_cont=5.1e-06 nfing=1 source_num=2 $X=-230840 $Y=-142980 $D=1
M11 4 6 4 4 nmos_a L=2e-06 W=0.0001 AD=7.86989e-13 AS=2.6e-11 PD=1.51344e-06 PS=1.51344e-06 w_cont=5.1e-06 nfing=1 source_num=2 $X=-220760 $Y=-142980 $D=1
M12 4 6 4 4 nmos_a L=2e-06 W=0.0001 AD=7.86989e-13 AS=2.6e-11 PD=1.51344e-06 PS=1.51344e-06 w_cont=5.1e-06 nfing=1 source_num=2 $X=-210680 $Y=-142980 $D=1
X14 4 6 ICV_146 $T=-308860 -143180 1 180 $X=-312060 $Y=-143180
X15 4 6 ICV_146 $T=-298780 -143180 1 180 $X=-301980 $Y=-143180
X16 4 6 ICV_146 $T=-288700 -143180 1 180 $X=-291900 $Y=-143180
X17 4 6 ICV_146 $T=-278620 -143180 1 180 $X=-281820 $Y=-143180
X18 4 6 ICV_146 $T=-268540 -143180 1 180 $X=-271740 $Y=-143180
X19 4 6 ICV_146 $T=-258460 -143180 1 180 $X=-261660 $Y=-143180
X20 4 6 ICV_146 $T=-248380 -143180 1 180 $X=-251580 $Y=-143180
X21 4 6 ICV_146 $T=-238300 -143180 1 180 $X=-241500 $Y=-143180
X22 4 6 ICV_146 $T=-228220 -143180 1 180 $X=-231420 $Y=-143180
X23 4 6 ICV_146 $T=-218140 -143180 1 180 $X=-221340 $Y=-143180
X24 4 6 ICV_146 $T=-208060 -143180 1 180 $X=-211260 $Y=-143180
.ENDS
***************************************
.SUBCKT ICV_156 2 4 5 6
** N=37 EP=4 IP=78 FDC=26
*.SEEDPROM
M0 20 20 21 21 nmos_a L=2.4e-07 W=1.2e-06 AD=7.2e-13 AS=4.8e-13 PD=1.8e-06 PS=9e-07 w_cont=6e-07 nfing=1 source_num=2 $X=-292400 $Y=-144820 $D=1
M1 22 22 6 6 nmos_a L=2.4e-07 W=1.2e-06 AD=7.2e-13 AS=4.8e-13 PD=1.8e-06 PS=9e-07 w_cont=6e-07 nfing=1 source_num=2 $X=-287000 $Y=-144820 $D=1
M2 23 23 24 24 nmos_a L=2.4e-07 W=1.2e-06 AD=7.2e-13 AS=4.8e-13 PD=1.8e-06 PS=9e-07 w_cont=6e-07 nfing=1 source_num=2 $X=-267200 $Y=-144820 $D=1
M3 25 25 6 6 nmos_a L=2.4e-07 W=1.2e-06 AD=7.2e-13 AS=4.8e-13 PD=1.8e-06 PS=9e-07 w_cont=6e-07 nfing=1 source_num=2 $X=-261800 $Y=-144820 $D=1
M4 26 26 27 27 nmos_a L=2.4e-07 W=1.2e-06 AD=7.2e-13 AS=4.8e-13 PD=1.8e-06 PS=9e-07 w_cont=6e-07 nfing=1 source_num=2 $X=-242000 $Y=-144820 $D=1
M5 28 28 6 6 nmos_a L=2.4e-07 W=1.2e-06 AD=7.2e-13 AS=4.8e-13 PD=1.8e-06 PS=9e-07 w_cont=6e-07 nfing=1 source_num=2 $X=-236600 $Y=-144820 $D=1
M6 29 29 30 30 nmos_a L=2.4e-07 W=1.2e-06 AD=7.2e-13 AS=4.8e-13 PD=1.8e-06 PS=9e-07 w_cont=6e-07 nfing=1 source_num=2 $X=-216800 $Y=-144820 $D=1
M7 31 31 6 6 nmos_a L=2.4e-07 W=1.2e-06 AD=7.2e-13 AS=4.8e-13 PD=1.8e-06 PS=9e-07 w_cont=6e-07 nfing=1 source_num=2 $X=-211400 $Y=-144820 $D=1
X8 5 4 5 pmos_a_CDNS_5887047866540 $T=-307360 -145440 0 90 $X=-309560 $Y=-145440
X9 5 20 20 pmos_a_CDNS_5887047866540 $T=-293100 -143960 1 270 $X=-295300 $Y=-145400
X10 21 22 22 pmos_a_CDNS_5887047866540 $T=-287700 -143960 1 270 $X=-289900 $Y=-145400
X11 5 4 5 pmos_a_CDNS_5887047866540 $T=-282160 -145440 0 90 $X=-284360 $Y=-145440
X12 5 23 23 pmos_a_CDNS_5887047866540 $T=-267900 -143960 1 270 $X=-270100 $Y=-145400
X13 24 25 25 pmos_a_CDNS_5887047866540 $T=-262500 -143960 1 270 $X=-264700 $Y=-145400
X14 5 4 5 pmos_a_CDNS_5887047866540 $T=-256960 -145440 0 90 $X=-259160 $Y=-145440
X15 5 26 26 pmos_a_CDNS_5887047866540 $T=-242700 -143960 1 270 $X=-244900 $Y=-145400
X16 27 28 28 pmos_a_CDNS_5887047866540 $T=-237300 -143960 1 270 $X=-239500 $Y=-145400
X17 5 4 5 pmos_a_CDNS_5887047866540 $T=-231760 -145440 0 90 $X=-233960 $Y=-145440
X18 5 29 29 pmos_a_CDNS_5887047866540 $T=-217500 -143960 1 270 $X=-219700 $Y=-145400
X19 30 31 31 pmos_a_CDNS_5887047866540 $T=-212100 -143960 1 270 $X=-214300 $Y=-145400
X20 5 4 5 pmos_a_CDNS_5887047866540 $T=-203500 -145440 0 90 $X=-205700 $Y=-145440
X29 4 2 5 nmos_a_CDNS_5887047866547 $T=-306780 -143960 0 270 $X=-306780 $Y=-145400
X30 4 2 5 nmos_a_CDNS_5887047866547 $T=-281580 -143960 0 270 $X=-281580 $Y=-145400
X31 4 2 5 nmos_a_CDNS_5887047866547 $T=-256380 -143960 0 270 $X=-256380 $Y=-145400
X32 4 2 5 nmos_a_CDNS_5887047866547 $T=-231180 -143960 0 270 $X=-231180 $Y=-145400
X33 4 2 5 nmos_a_CDNS_5887047866547 $T=-202920 -143960 0 270 $X=-202920 $Y=-145400
.ENDS
***************************************
.SUBCKT ICV_157 1 2 3 4
** N=4 EP=4 IP=8 FDC=22
*.SEEDPROM
M0 1 4 4 4 pmos_a L=2.4e-07 W=1e-06 AD=5.928e-13 AS=1.61e-13 PD=1.6e-06 PS=8e-07 w_cont=6e-07 nfing=1 mmm=1 $X=11580 $Y=-1960 $D=5
M1 1 4 4 4 pmos_a L=2.4e-07 W=1e-06 AD=5.928e-13 AS=1.61e-13 PD=1.6e-06 PS=8e-07 w_cont=6e-07 nfing=1 mmm=1 $X=11580 $Y=360 $D=5
X2 1 2 3 4 ICV_149 $T=0 0 1 0 $X=-360 $Y=-3220
X3 1 2 3 4 ICV_149 $T=0 0 0 0 $X=-360 $Y=-340
.ENDS
***************************************
.SUBCKT ICV_158 1 2 3 4
** N=4 EP=4 IP=8 FDC=46
*.SEEDPROM
M0 3 4 4 4 pmos_a L=2.4e-07 W=1e-06 AD=5.928e-13 AS=1.61e-13 PD=1.6e-06 PS=8e-07 w_cont=6e-07 nfing=1 mmm=1 $X=12340 $Y=-1960 $D=5
M1 3 4 4 4 pmos_a L=2.4e-07 W=1e-06 AD=5.928e-13 AS=1.61e-13 PD=1.6e-06 PS=8e-07 w_cont=6e-07 nfing=1 mmm=1 $X=12340 $Y=360 $D=5
X2 3 2 1 4 ICV_157 $T=0 0 0 0 $X=-360 $Y=-3220
X3 3 2 1 4 ICV_157 $T=12080 0 0 0 $X=11720 $Y=-3220
.ENDS
***************************************
.SUBCKT ICV_159 1 2 3 4
** N=4 EP=4 IP=8 FDC=94
*.SEEDPROM
M0 3 4 4 4 pmos_a L=2.4e-07 W=1e-06 AD=5.928e-13 AS=1.61e-13 PD=1.6e-06 PS=8e-07 w_cont=6e-07 nfing=1 mmm=1 $X=24420 $Y=-1960 $D=5
M1 3 4 4 4 pmos_a L=2.4e-07 W=1e-06 AD=5.928e-13 AS=1.61e-13 PD=1.6e-06 PS=8e-07 w_cont=6e-07 nfing=1 mmm=1 $X=24420 $Y=360 $D=5
X2 1 2 3 4 ICV_158 $T=0 0 0 0 $X=-360 $Y=-3220
X3 1 2 3 4 ICV_158 $T=24160 0 0 0 $X=23800 $Y=-3220
.ENDS
***************************************
.SUBCKT ICV_160 1 2 3 13 14 15 16 17
** N=18 EP=8 IP=66 FDC=1706
*.SEEDPROM
M0 18 1 2 2 nmos_a L=2.8e-07 W=4.8e-07 AD=4.32e-13 AS=1.92e-13 PD=1.08e-06 PS=5.4e-07 w_cont=6e-07 nfing=1 source_num=2 $X=-1010020 $Y=270000 $D=1
M1 13 13 2 2 nmos_a L=2.4e-07 W=4.8e-07 AD=4.32e-13 AS=1.92e-13 PD=1.08e-06 PS=5.4e-07 w_cont=6e-07 nfing=1 source_num=2 $X=-1008800 $Y=268500 $D=1
M2 15 18 14 14 nmos_a L=2.8e-07 W=4.8e-07 AD=4.32e-13 AS=1.92e-13 PD=1.08e-06 PS=5.4e-07 w_cont=6e-07 nfing=1 source_num=2 $X=-1008540 $Y=271480 $D=1
M3 14 16 2 2 nmos_a L=2.4e-07 W=1.2e-06 AD=7.2e-13 AS=4.8e-13 PD=1.8e-06 PS=9e-07 w_cont=6e-07 nfing=1 source_num=2 $X=-1008800 $Y=273600 $D=1
M4 18 1 3 3 pmos_a L=2.8e-07 W=4.8e-07 AD=4.32e-13 AS=1.224e-13 PD=1.08e-06 PS=5.4e-07 w_cont=6e-07 nfing=1 mmm=1 $X=-1010020 $Y=271980 $D=5
M5 17 16 16 16 pmos_a L=2.4e-07 W=1e-06 AD=5.928e-13 AS=1.61e-13 PD=1.6e-06 PS=8e-07 w_cont=6e-07 nfing=1 mmm=1 $X=-401620 $Y=269800 $D=5
M6 17 16 16 16 pmos_a L=2.4e-07 W=1e-06 AD=5.928e-13 AS=1.61e-13 PD=1.6e-06 PS=8e-07 w_cont=6e-07 nfing=1 mmm=1 $X=-396340 $Y=269800 $D=5
M7 17 16 16 16 pmos_a L=2.4e-07 W=1e-06 AD=5.928e-13 AS=1.61e-13 PD=1.6e-06 PS=8e-07 w_cont=6e-07 nfing=1 mmm=1 $X=-401620 $Y=272120 $D=5
M8 17 16 16 16 pmos_a L=2.4e-07 W=1e-06 AD=5.928e-13 AS=1.61e-13 PD=1.6e-06 PS=8e-07 w_cont=6e-07 nfing=1 mmm=1 $X=-396340 $Y=272120 $D=5
M9 17 16 16 16 pmos_a L=2.4e-07 W=1e-06 AD=5.928e-13 AS=1.61e-13 PD=1.6e-06 PS=8e-07 w_cont=6e-07 nfing=1 mmm=1 $X=-425780 $Y=272120 $D=5
M10 17 16 16 16 pmos_a L=2.4e-07 W=1e-06 AD=5.928e-13 AS=1.61e-13 PD=1.6e-06 PS=8e-07 w_cont=6e-07 nfing=1 mmm=1 $X=-425780 $Y=269800 $D=5
M11 17 16 16 16 pmos_a L=2.4e-07 W=1e-06 AD=5.928e-13 AS=1.25e-13 PD=1.6e-06 PS=8e-07 w_cont=6e-07 nfing=1 mmm=1 $X=-1005620 $Y=272120 $D=5
M12 17 16 16 16 pmos_a L=2.4e-07 W=1e-06 AD=5.928e-13 AS=1.25e-13 PD=1.6e-06 PS=8e-07 w_cont=6e-07 nfing=1 mmm=1 $X=-1005620 $Y=269800 $D=5
M13 17 16 16 16 pmos_a L=2.4e-07 W=1e-06 AD=5.928e-13 AS=1.61e-13 PD=1.6e-06 PS=8e-07 w_cont=6e-07 nfing=1 mmm=1 $X=-957300 $Y=272120 $D=5
M14 17 16 16 16 pmos_a L=2.4e-07 W=1e-06 AD=5.928e-13 AS=1.61e-13 PD=1.6e-06 PS=8e-07 w_cont=6e-07 nfing=1 mmm=1 $X=-957300 $Y=269800 $D=5
M15 17 16 16 16 pmos_a L=2.4e-07 W=1e-06 AD=5.928e-13 AS=1.61e-13 PD=1.6e-06 PS=8e-07 w_cont=6e-07 nfing=1 mmm=1 $X=-908980 $Y=272120 $D=5
M16 17 16 16 16 pmos_a L=2.4e-07 W=1e-06 AD=5.928e-13 AS=1.61e-13 PD=1.6e-06 PS=8e-07 w_cont=6e-07 nfing=1 mmm=1 $X=-908980 $Y=269800 $D=5
M17 17 16 16 16 pmos_a L=2.4e-07 W=1e-06 AD=5.928e-13 AS=1.61e-13 PD=1.6e-06 PS=8e-07 w_cont=6e-07 nfing=1 mmm=1 $X=-860660 $Y=272120 $D=5
M18 17 16 16 16 pmos_a L=2.4e-07 W=1e-06 AD=5.928e-13 AS=1.61e-13 PD=1.6e-06 PS=8e-07 w_cont=6e-07 nfing=1 mmm=1 $X=-860660 $Y=269800 $D=5
M19 17 16 16 16 pmos_a L=2.4e-07 W=1e-06 AD=5.928e-13 AS=1.61e-13 PD=1.6e-06 PS=8e-07 w_cont=6e-07 nfing=1 mmm=1 $X=-812340 $Y=272120 $D=5
M20 17 16 16 16 pmos_a L=2.4e-07 W=1e-06 AD=5.928e-13 AS=1.61e-13 PD=1.6e-06 PS=8e-07 w_cont=6e-07 nfing=1 mmm=1 $X=-812340 $Y=269800 $D=5
M21 17 16 16 16 pmos_a L=2.4e-07 W=1e-06 AD=5.928e-13 AS=1.61e-13 PD=1.6e-06 PS=8e-07 w_cont=6e-07 nfing=1 mmm=1 $X=-764020 $Y=272120 $D=5
M22 17 16 16 16 pmos_a L=2.4e-07 W=1e-06 AD=5.928e-13 AS=1.61e-13 PD=1.6e-06 PS=8e-07 w_cont=6e-07 nfing=1 mmm=1 $X=-764020 $Y=269800 $D=5
M23 17 16 16 16 pmos_a L=2.4e-07 W=1e-06 AD=5.928e-13 AS=1.61e-13 PD=1.6e-06 PS=8e-07 w_cont=6e-07 nfing=1 mmm=1 $X=-715700 $Y=272120 $D=5
M24 17 16 16 16 pmos_a L=2.4e-07 W=1e-06 AD=5.928e-13 AS=1.61e-13 PD=1.6e-06 PS=8e-07 w_cont=6e-07 nfing=1 mmm=1 $X=-715700 $Y=269800 $D=5
M25 17 16 16 16 pmos_a L=2.4e-07 W=1e-06 AD=5.928e-13 AS=1.61e-13 PD=1.6e-06 PS=8e-07 w_cont=6e-07 nfing=1 mmm=1 $X=-667380 $Y=272120 $D=5
M26 17 16 16 16 pmos_a L=2.4e-07 W=1e-06 AD=5.928e-13 AS=1.61e-13 PD=1.6e-06 PS=8e-07 w_cont=6e-07 nfing=1 mmm=1 $X=-667380 $Y=269800 $D=5
M27 17 16 16 16 pmos_a L=2.4e-07 W=1e-06 AD=5.928e-13 AS=1.61e-13 PD=1.6e-06 PS=8e-07 w_cont=6e-07 nfing=1 mmm=1 $X=-619060 $Y=272120 $D=5
M28 17 16 16 16 pmos_a L=2.4e-07 W=1e-06 AD=5.928e-13 AS=1.61e-13 PD=1.6e-06 PS=8e-07 w_cont=6e-07 nfing=1 mmm=1 $X=-619060 $Y=269800 $D=5
M29 17 16 16 16 pmos_a L=2.4e-07 W=1e-06 AD=5.928e-13 AS=1.61e-13 PD=1.6e-06 PS=8e-07 w_cont=6e-07 nfing=1 mmm=1 $X=-570740 $Y=272120 $D=5
M30 17 16 16 16 pmos_a L=2.4e-07 W=1e-06 AD=5.928e-13 AS=1.61e-13 PD=1.6e-06 PS=8e-07 w_cont=6e-07 nfing=1 mmm=1 $X=-570740 $Y=269800 $D=5
M31 17 16 16 16 pmos_a L=2.4e-07 W=1e-06 AD=5.928e-13 AS=1.61e-13 PD=1.6e-06 PS=8e-07 w_cont=6e-07 nfing=1 mmm=1 $X=-522420 $Y=272120 $D=5
M32 17 16 16 16 pmos_a L=2.4e-07 W=1e-06 AD=5.928e-13 AS=1.61e-13 PD=1.6e-06 PS=8e-07 w_cont=6e-07 nfing=1 mmm=1 $X=-522420 $Y=269800 $D=5
M33 17 16 16 16 pmos_a L=2.4e-07 W=1e-06 AD=5.928e-13 AS=1.61e-13 PD=1.6e-06 PS=8e-07 w_cont=6e-07 nfing=1 mmm=1 $X=-474100 $Y=272120 $D=5
M34 17 16 16 16 pmos_a L=2.4e-07 W=1e-06 AD=5.928e-13 AS=1.61e-13 PD=1.6e-06 PS=8e-07 w_cont=6e-07 nfing=1 mmm=1 $X=-474100 $Y=269800 $D=5
M35 2 3 2 cpoly_p w=3.8e-06 l=2e-06 c=5.2038e-14 as=1.81137e-13 ad=7.488e-13 ps=1.44e-06 pd=1.11673e-06 sim_w=2.88e-06 m_per_maxw=1.31944 numb_sub_cont=3 nfing=1 $X=-1013500 $Y=276580 $D=21
M36 2 3 2 cpoly_p w=3.8e-06 l=2e-06 c=5.2038e-14 as=2.31158e-13 ad=7.488e-13 ps=1.44e-06 pd=1.11673e-06 sim_w=2.88e-06 m_per_maxw=1.31944 numb_sub_cont=3 nfing=1 $X=-1010980 $Y=276580 $D=21
M37 2 3 2 cpoly_p w=3.8e-06 l=2e-06 c=5.2038e-14 as=2.31158e-13 ad=7.488e-13 ps=1.44e-06 pd=1.11673e-06 sim_w=2.88e-06 m_per_maxw=1.31944 numb_sub_cont=3 nfing=1 $X=-1008460 $Y=276580 $D=21
M38 2 3 2 cpoly_p w=3.8e-06 l=2e-06 c=5.2038e-14 as=2.31158e-13 ad=7.488e-13 ps=1.44e-06 pd=1.11673e-06 sim_w=2.88e-06 m_per_maxw=1.31944 numb_sub_cont=3 nfing=1 $X=-1005940 $Y=276580 $D=21
M39 2 3 2 cpoly_p w=3.8e-06 l=2e-06 c=5.2038e-14 as=2.31158e-13 ad=7.488e-13 ps=1.44e-06 pd=1.11673e-06 sim_w=2.88e-06 m_per_maxw=1.31944 numb_sub_cont=3 nfing=1 $X=-1003420 $Y=276580 $D=21
M40 2 3 2 cpoly_p w=3.8e-06 l=2e-06 c=5.2038e-14 as=2.31158e-13 ad=7.488e-13 ps=1.44e-06 pd=1.11673e-06 sim_w=2.88e-06 m_per_maxw=1.31944 numb_sub_cont=3 nfing=1 $X=-1000900 $Y=276580 $D=21
M41 2 3 2 cpoly_p w=3.8e-06 l=2e-06 c=5.2038e-14 as=2.31158e-13 ad=7.488e-13 ps=1.44e-06 pd=1.11673e-06 sim_w=2.88e-06 m_per_maxw=1.31944 numb_sub_cont=3 nfing=1 $X=-998380 $Y=276580 $D=21
M42 2 3 2 cpoly_p w=3.8e-06 l=2e-06 c=5.2038e-14 as=2.31158e-13 ad=7.488e-13 ps=1.44e-06 pd=1.11673e-06 sim_w=2.88e-06 m_per_maxw=1.31944 numb_sub_cont=3 nfing=1 $X=-995860 $Y=276580 $D=21
M43 2 3 2 cpoly_p w=3.8e-06 l=2e-06 c=5.2038e-14 as=2.31158e-13 ad=7.488e-13 ps=1.44e-06 pd=1.11673e-06 sim_w=2.88e-06 m_per_maxw=1.31944 numb_sub_cont=3 nfing=1 $X=-993340 $Y=276580 $D=21
M44 2 3 2 cpoly_p w=3.8e-06 l=2e-06 c=5.2038e-14 as=2.31158e-13 ad=7.488e-13 ps=1.44e-06 pd=1.11673e-06 sim_w=2.88e-06 m_per_maxw=1.31944 numb_sub_cont=3 nfing=1 $X=-990820 $Y=276580 $D=21
M45 2 3 2 cpoly_p w=3.8e-06 l=2e-06 c=5.2038e-14 as=2.31158e-13 ad=7.488e-13 ps=1.44e-06 pd=1.11673e-06 sim_w=2.88e-06 m_per_maxw=1.31944 numb_sub_cont=3 nfing=1 $X=-988300 $Y=276580 $D=21
M46 2 3 2 cpoly_p w=3.8e-06 l=2e-06 c=5.2038e-14 as=2.31158e-13 ad=7.488e-13 ps=1.44e-06 pd=1.11673e-06 sim_w=2.88e-06 m_per_maxw=1.31944 numb_sub_cont=3 nfing=1 $X=-985780 $Y=276580 $D=21
M47 2 3 2 cpoly_p w=3.8e-06 l=2e-06 c=5.2038e-14 as=2.31158e-13 ad=7.488e-13 ps=1.44e-06 pd=1.11673e-06 sim_w=2.88e-06 m_per_maxw=1.31944 numb_sub_cont=3 nfing=1 $X=-983260 $Y=276580 $D=21
M48 2 3 2 cpoly_p w=3.8e-06 l=2e-06 c=5.2038e-14 as=2.31158e-13 ad=7.488e-13 ps=1.44e-06 pd=1.11673e-06 sim_w=2.88e-06 m_per_maxw=1.31944 numb_sub_cont=3 nfing=1 $X=-980740 $Y=276580 $D=21
M49 2 3 2 cpoly_p w=3.8e-06 l=2e-06 c=5.2038e-14 as=2.31158e-13 ad=7.488e-13 ps=1.44e-06 pd=1.11673e-06 sim_w=2.88e-06 m_per_maxw=1.31944 numb_sub_cont=3 nfing=1 $X=-978220 $Y=276580 $D=21
M50 2 3 2 cpoly_p w=3.8e-06 l=2e-06 c=5.2038e-14 as=2.31158e-13 ad=7.488e-13 ps=1.44e-06 pd=1.11673e-06 sim_w=2.88e-06 m_per_maxw=1.31944 numb_sub_cont=3 nfing=1 $X=-975700 $Y=276580 $D=21
M51 2 3 2 cpoly_p w=3.8e-06 l=2e-06 c=5.2038e-14 as=2.31158e-13 ad=7.488e-13 ps=1.44e-06 pd=1.11673e-06 sim_w=2.88e-06 m_per_maxw=1.31944 numb_sub_cont=3 nfing=1 $X=-973180 $Y=276580 $D=21
M52 2 3 2 cpoly_p w=3.8e-06 l=2e-06 c=5.2038e-14 as=2.31158e-13 ad=7.488e-13 ps=1.44e-06 pd=1.11673e-06 sim_w=2.88e-06 m_per_maxw=1.31944 numb_sub_cont=3 nfing=1 $X=-970660 $Y=276580 $D=21
M53 2 3 2 cpoly_p w=3.8e-06 l=2e-06 c=5.2038e-14 as=2.31158e-13 ad=7.488e-13 ps=1.44e-06 pd=1.11673e-06 sim_w=2.88e-06 m_per_maxw=1.31944 numb_sub_cont=3 nfing=1 $X=-968140 $Y=276580 $D=21
M54 2 3 2 cpoly_p w=3.8e-06 l=2e-06 c=5.2038e-14 as=2.31158e-13 ad=7.488e-13 ps=1.44e-06 pd=1.11673e-06 sim_w=2.88e-06 m_per_maxw=1.31944 numb_sub_cont=3 nfing=1 $X=-965620 $Y=276580 $D=21
M55 2 3 2 cpoly_p w=3.8e-06 l=2e-06 c=5.2038e-14 as=2.31158e-13 ad=7.488e-13 ps=1.44e-06 pd=1.11673e-06 sim_w=2.88e-06 m_per_maxw=1.31944 numb_sub_cont=3 nfing=1 $X=-963100 $Y=276580 $D=21
M56 2 3 2 cpoly_p w=3.8e-06 l=2e-06 c=5.2038e-14 as=2.31158e-13 ad=7.488e-13 ps=1.44e-06 pd=1.11673e-06 sim_w=2.88e-06 m_per_maxw=1.31944 numb_sub_cont=3 nfing=1 $X=-960580 $Y=276580 $D=21
M57 2 3 2 cpoly_p w=3.8e-06 l=2e-06 c=5.2038e-14 as=2.31158e-13 ad=7.488e-13 ps=1.44e-06 pd=1.11673e-06 sim_w=2.88e-06 m_per_maxw=1.31944 numb_sub_cont=3 nfing=1 $X=-958060 $Y=276580 $D=21
M58 2 3 2 cpoly_p w=3.8e-06 l=2e-06 c=5.2038e-14 as=2.31158e-13 ad=7.488e-13 ps=1.44e-06 pd=1.11673e-06 sim_w=2.88e-06 m_per_maxw=1.31944 numb_sub_cont=3 nfing=1 $X=-955540 $Y=276580 $D=21
M59 2 3 2 cpoly_p w=3.8e-06 l=2e-06 c=5.2038e-14 as=2.31158e-13 ad=7.488e-13 ps=1.44e-06 pd=1.11673e-06 sim_w=2.88e-06 m_per_maxw=1.31944 numb_sub_cont=3 nfing=1 $X=-953020 $Y=276580 $D=21
M60 2 3 2 cpoly_p w=3.8e-06 l=2e-06 c=5.2038e-14 as=2.31158e-13 ad=7.488e-13 ps=1.44e-06 pd=1.11673e-06 sim_w=2.88e-06 m_per_maxw=1.31944 numb_sub_cont=3 nfing=1 $X=-950500 $Y=276580 $D=21
M61 2 3 2 cpoly_p w=3.8e-06 l=2e-06 c=5.2038e-14 as=2.31158e-13 ad=7.488e-13 ps=1.44e-06 pd=1.11673e-06 sim_w=2.88e-06 m_per_maxw=1.31944 numb_sub_cont=3 nfing=1 $X=-947980 $Y=276580 $D=21
M62 2 3 2 cpoly_p w=3.8e-06 l=2e-06 c=5.2038e-14 as=2.31158e-13 ad=7.488e-13 ps=1.44e-06 pd=1.11673e-06 sim_w=2.88e-06 m_per_maxw=1.31944 numb_sub_cont=3 nfing=1 $X=-945460 $Y=276580 $D=21
M63 2 3 2 cpoly_p w=3.8e-06 l=2e-06 c=5.2038e-14 as=2.31158e-13 ad=7.488e-13 ps=1.44e-06 pd=1.11673e-06 sim_w=2.88e-06 m_per_maxw=1.31944 numb_sub_cont=3 nfing=1 $X=-942940 $Y=276580 $D=21
M64 2 3 2 cpoly_p w=3.8e-06 l=2e-06 c=5.2038e-14 as=2.31158e-13 ad=7.488e-13 ps=1.44e-06 pd=1.11673e-06 sim_w=2.88e-06 m_per_maxw=1.31944 numb_sub_cont=3 nfing=1 $X=-940420 $Y=276580 $D=21
M65 2 3 2 cpoly_p w=3.8e-06 l=2e-06 c=5.2038e-14 as=2.31158e-13 ad=7.488e-13 ps=1.44e-06 pd=1.11673e-06 sim_w=2.88e-06 m_per_maxw=1.31944 numb_sub_cont=3 nfing=1 $X=-937900 $Y=276580 $D=21
M66 2 3 2 cpoly_p w=3.8e-06 l=2e-06 c=5.2038e-14 as=2.31158e-13 ad=7.488e-13 ps=1.44e-06 pd=1.11673e-06 sim_w=2.88e-06 m_per_maxw=1.31944 numb_sub_cont=3 nfing=1 $X=-935380 $Y=276580 $D=21
M67 2 3 2 cpoly_p w=3.8e-06 l=2e-06 c=5.2038e-14 as=2.31158e-13 ad=7.488e-13 ps=1.44e-06 pd=1.11673e-06 sim_w=2.88e-06 m_per_maxw=1.31944 numb_sub_cont=3 nfing=1 $X=-932860 $Y=276580 $D=21
M68 2 3 2 cpoly_p w=3.8e-06 l=2e-06 c=5.2038e-14 as=2.31158e-13 ad=7.488e-13 ps=1.44e-06 pd=1.11673e-06 sim_w=2.88e-06 m_per_maxw=1.31944 numb_sub_cont=3 nfing=1 $X=-930340 $Y=276580 $D=21
M69 2 3 2 cpoly_p w=3.8e-06 l=2e-06 c=5.2038e-14 as=2.31158e-13 ad=7.488e-13 ps=1.44e-06 pd=1.11673e-06 sim_w=2.88e-06 m_per_maxw=1.31944 numb_sub_cont=3 nfing=1 $X=-927820 $Y=276580 $D=21
M70 2 3 2 cpoly_p w=3.8e-06 l=2e-06 c=5.2038e-14 as=2.31158e-13 ad=7.488e-13 ps=1.44e-06 pd=1.11673e-06 sim_w=2.88e-06 m_per_maxw=1.31944 numb_sub_cont=3 nfing=1 $X=-925300 $Y=276580 $D=21
M71 2 3 2 cpoly_p w=3.8e-06 l=2e-06 c=5.2038e-14 as=2.31158e-13 ad=7.488e-13 ps=1.44e-06 pd=1.11673e-06 sim_w=2.88e-06 m_per_maxw=1.31944 numb_sub_cont=3 nfing=1 $X=-922780 $Y=276580 $D=21
M72 2 3 2 cpoly_p w=3.8e-06 l=2e-06 c=5.2038e-14 as=2.31158e-13 ad=7.488e-13 ps=1.44e-06 pd=1.11673e-06 sim_w=2.88e-06 m_per_maxw=1.31944 numb_sub_cont=3 nfing=1 $X=-920260 $Y=276580 $D=21
M73 2 3 2 cpoly_p w=3.8e-06 l=2e-06 c=5.2038e-14 as=2.31158e-13 ad=7.488e-13 ps=1.44e-06 pd=1.11673e-06 sim_w=2.88e-06 m_per_maxw=1.31944 numb_sub_cont=3 nfing=1 $X=-917740 $Y=276580 $D=21
M74 2 3 2 cpoly_p w=3.8e-06 l=2e-06 c=5.2038e-14 as=2.31158e-13 ad=7.488e-13 ps=1.44e-06 pd=1.11673e-06 sim_w=2.88e-06 m_per_maxw=1.31944 numb_sub_cont=3 nfing=1 $X=-915220 $Y=276580 $D=21
M75 2 3 2 cpoly_p w=3.8e-06 l=2e-06 c=5.2038e-14 as=2.31158e-13 ad=7.488e-13 ps=1.44e-06 pd=1.11673e-06 sim_w=2.88e-06 m_per_maxw=1.31944 numb_sub_cont=3 nfing=1 $X=-912700 $Y=276580 $D=21
M76 2 3 2 cpoly_p w=3.8e-06 l=2e-06 c=5.2038e-14 as=2.31158e-13 ad=7.488e-13 ps=1.44e-06 pd=1.11673e-06 sim_w=2.88e-06 m_per_maxw=1.31944 numb_sub_cont=3 nfing=1 $X=-910180 $Y=276580 $D=21
M77 2 3 2 cpoly_p w=3.8e-06 l=2e-06 c=5.2038e-14 as=2.31158e-13 ad=7.488e-13 ps=1.44e-06 pd=1.11673e-06 sim_w=2.88e-06 m_per_maxw=1.31944 numb_sub_cont=3 nfing=1 $X=-907660 $Y=276580 $D=21
M78 2 3 2 cpoly_p w=3.8e-06 l=2e-06 c=5.2038e-14 as=2.31158e-13 ad=7.488e-13 ps=1.44e-06 pd=1.11673e-06 sim_w=2.88e-06 m_per_maxw=1.31944 numb_sub_cont=3 nfing=1 $X=-905140 $Y=276580 $D=21
M79 2 3 2 cpoly_p w=3.8e-06 l=2e-06 c=5.2038e-14 as=2.31158e-13 ad=7.488e-13 ps=1.44e-06 pd=1.11673e-06 sim_w=2.88e-06 m_per_maxw=1.31944 numb_sub_cont=3 nfing=1 $X=-902620 $Y=276580 $D=21
M80 2 3 2 cpoly_p w=3.8e-06 l=2e-06 c=5.2038e-14 as=2.31158e-13 ad=7.488e-13 ps=1.44e-06 pd=1.11673e-06 sim_w=2.88e-06 m_per_maxw=1.31944 numb_sub_cont=3 nfing=1 $X=-900100 $Y=276580 $D=21
M81 2 3 2 cpoly_p w=3.8e-06 l=2e-06 c=5.2038e-14 as=2.31158e-13 ad=7.488e-13 ps=1.44e-06 pd=1.11673e-06 sim_w=2.88e-06 m_per_maxw=1.31944 numb_sub_cont=3 nfing=1 $X=-897580 $Y=276580 $D=21
M82 2 3 2 cpoly_p w=3.8e-06 l=2e-06 c=5.2038e-14 as=2.31158e-13 ad=7.488e-13 ps=1.44e-06 pd=1.11673e-06 sim_w=2.88e-06 m_per_maxw=1.31944 numb_sub_cont=3 nfing=1 $X=-895060 $Y=276580 $D=21
M83 2 3 2 cpoly_p w=3.8e-06 l=2e-06 c=5.2038e-14 as=2.31158e-13 ad=7.488e-13 ps=1.44e-06 pd=1.11673e-06 sim_w=2.88e-06 m_per_maxw=1.31944 numb_sub_cont=3 nfing=1 $X=-892540 $Y=276580 $D=21
M84 2 3 2 cpoly_p w=3.8e-06 l=2e-06 c=5.2038e-14 as=2.31158e-13 ad=7.488e-13 ps=1.44e-06 pd=1.11673e-06 sim_w=2.88e-06 m_per_maxw=1.31944 numb_sub_cont=3 nfing=1 $X=-890020 $Y=276580 $D=21
M85 2 3 2 cpoly_p w=3.8e-06 l=2e-06 c=5.2038e-14 as=2.31158e-13 ad=7.488e-13 ps=1.44e-06 pd=1.11673e-06 sim_w=2.88e-06 m_per_maxw=1.31944 numb_sub_cont=3 nfing=1 $X=-887500 $Y=276580 $D=21
M86 2 3 2 cpoly_p w=3.8e-06 l=2e-06 c=5.2038e-14 as=2.31158e-13 ad=7.488e-13 ps=1.44e-06 pd=1.11673e-06 sim_w=2.88e-06 m_per_maxw=1.31944 numb_sub_cont=3 nfing=1 $X=-884980 $Y=276580 $D=21
M87 2 3 2 cpoly_p w=3.8e-06 l=2e-06 c=5.2038e-14 as=2.31158e-13 ad=7.488e-13 ps=1.44e-06 pd=1.11673e-06 sim_w=2.88e-06 m_per_maxw=1.31944 numb_sub_cont=3 nfing=1 $X=-882460 $Y=276580 $D=21
M88 2 3 2 cpoly_p w=3.8e-06 l=2e-06 c=5.2038e-14 as=2.31158e-13 ad=7.488e-13 ps=1.44e-06 pd=1.11673e-06 sim_w=2.88e-06 m_per_maxw=1.31944 numb_sub_cont=3 nfing=1 $X=-879940 $Y=276580 $D=21
M89 2 3 2 cpoly_p w=3.8e-06 l=2e-06 c=5.2038e-14 as=2.31158e-13 ad=7.488e-13 ps=1.44e-06 pd=1.11673e-06 sim_w=2.88e-06 m_per_maxw=1.31944 numb_sub_cont=3 nfing=1 $X=-877420 $Y=276580 $D=21
M90 2 3 2 cpoly_p w=3.8e-06 l=2e-06 c=5.2038e-14 as=2.31158e-13 ad=7.488e-13 ps=1.44e-06 pd=1.11673e-06 sim_w=2.88e-06 m_per_maxw=1.31944 numb_sub_cont=3 nfing=1 $X=-874900 $Y=276580 $D=21
M91 2 3 2 cpoly_p w=3.8e-06 l=2e-06 c=5.2038e-14 as=2.31158e-13 ad=7.488e-13 ps=1.44e-06 pd=1.11673e-06 sim_w=2.88e-06 m_per_maxw=1.31944 numb_sub_cont=3 nfing=1 $X=-872380 $Y=276580 $D=21
M92 2 3 2 cpoly_p w=3.8e-06 l=2e-06 c=5.2038e-14 as=2.31158e-13 ad=7.488e-13 ps=1.44e-06 pd=1.11673e-06 sim_w=2.88e-06 m_per_maxw=1.31944 numb_sub_cont=3 nfing=1 $X=-869860 $Y=276580 $D=21
M93 2 3 2 cpoly_p w=3.8e-06 l=2e-06 c=5.2038e-14 as=2.31158e-13 ad=7.488e-13 ps=1.44e-06 pd=1.11673e-06 sim_w=2.88e-06 m_per_maxw=1.31944 numb_sub_cont=3 nfing=1 $X=-867340 $Y=276580 $D=21
M94 2 3 2 cpoly_p w=3.8e-06 l=2e-06 c=5.2038e-14 as=2.31158e-13 ad=7.488e-13 ps=1.44e-06 pd=1.11673e-06 sim_w=2.88e-06 m_per_maxw=1.31944 numb_sub_cont=3 nfing=1 $X=-864820 $Y=276580 $D=21
M95 2 3 2 cpoly_p w=3.8e-06 l=2e-06 c=5.2038e-14 as=2.31158e-13 ad=7.488e-13 ps=1.44e-06 pd=1.11673e-06 sim_w=2.88e-06 m_per_maxw=1.31944 numb_sub_cont=3 nfing=1 $X=-862300 $Y=276580 $D=21
M96 2 3 2 cpoly_p w=3.8e-06 l=2e-06 c=5.2038e-14 as=2.31158e-13 ad=7.488e-13 ps=1.44e-06 pd=1.11673e-06 sim_w=2.88e-06 m_per_maxw=1.31944 numb_sub_cont=3 nfing=1 $X=-859780 $Y=276580 $D=21
M97 2 3 2 cpoly_p w=3.8e-06 l=2e-06 c=5.2038e-14 as=2.31158e-13 ad=7.488e-13 ps=1.44e-06 pd=1.11673e-06 sim_w=2.88e-06 m_per_maxw=1.31944 numb_sub_cont=3 nfing=1 $X=-857260 $Y=276580 $D=21
M98 2 3 2 cpoly_p w=3.8e-06 l=2e-06 c=5.2038e-14 as=2.31158e-13 ad=7.488e-13 ps=1.44e-06 pd=1.11673e-06 sim_w=2.88e-06 m_per_maxw=1.31944 numb_sub_cont=3 nfing=1 $X=-854740 $Y=276580 $D=21
M99 2 3 2 cpoly_p w=3.8e-06 l=2e-06 c=5.2038e-14 as=2.31158e-13 ad=7.488e-13 ps=1.44e-06 pd=1.11673e-06 sim_w=2.88e-06 m_per_maxw=1.31944 numb_sub_cont=3 nfing=1 $X=-852220 $Y=276580 $D=21
M100 2 3 2 cpoly_p w=3.8e-06 l=2e-06 c=5.2038e-14 as=2.31158e-13 ad=7.488e-13 ps=1.44e-06 pd=1.11673e-06 sim_w=2.88e-06 m_per_maxw=1.31944 numb_sub_cont=3 nfing=1 $X=-849700 $Y=276580 $D=21
M101 2 3 2 cpoly_p w=3.8e-06 l=2e-06 c=5.2038e-14 as=2.31158e-13 ad=7.488e-13 ps=1.44e-06 pd=1.11673e-06 sim_w=2.88e-06 m_per_maxw=1.31944 numb_sub_cont=3 nfing=1 $X=-847180 $Y=276580 $D=21
M102 2 3 2 cpoly_p w=3.8e-06 l=2e-06 c=5.2038e-14 as=2.31158e-13 ad=7.488e-13 ps=1.44e-06 pd=1.11673e-06 sim_w=2.88e-06 m_per_maxw=1.31944 numb_sub_cont=3 nfing=1 $X=-844660 $Y=276580 $D=21
M103 2 3 2 cpoly_p w=3.8e-06 l=2e-06 c=5.2038e-14 as=2.31158e-13 ad=7.488e-13 ps=1.44e-06 pd=1.11673e-06 sim_w=2.88e-06 m_per_maxw=1.31944 numb_sub_cont=3 nfing=1 $X=-842140 $Y=276580 $D=21
M104 2 3 2 cpoly_p w=3.8e-06 l=2e-06 c=5.2038e-14 as=2.31158e-13 ad=7.488e-13 ps=1.44e-06 pd=1.11673e-06 sim_w=2.88e-06 m_per_maxw=1.31944 numb_sub_cont=3 nfing=1 $X=-839620 $Y=276580 $D=21
M105 2 3 2 cpoly_p w=3.8e-06 l=2e-06 c=5.2038e-14 as=2.31158e-13 ad=7.488e-13 ps=1.44e-06 pd=1.11673e-06 sim_w=2.88e-06 m_per_maxw=1.31944 numb_sub_cont=3 nfing=1 $X=-837100 $Y=276580 $D=21
M106 2 3 2 cpoly_p w=3.8e-06 l=2e-06 c=5.2038e-14 as=2.31158e-13 ad=7.488e-13 ps=1.44e-06 pd=1.11673e-06 sim_w=2.88e-06 m_per_maxw=1.31944 numb_sub_cont=3 nfing=1 $X=-834580 $Y=276580 $D=21
M107 2 3 2 cpoly_p w=3.8e-06 l=2e-06 c=5.2038e-14 as=2.31158e-13 ad=7.488e-13 ps=1.44e-06 pd=1.11673e-06 sim_w=2.88e-06 m_per_maxw=1.31944 numb_sub_cont=3 nfing=1 $X=-832060 $Y=276580 $D=21
M108 2 3 2 cpoly_p w=3.8e-06 l=2e-06 c=5.2038e-14 as=2.31158e-13 ad=7.488e-13 ps=1.44e-06 pd=1.11673e-06 sim_w=2.88e-06 m_per_maxw=1.31944 numb_sub_cont=3 nfing=1 $X=-829540 $Y=276580 $D=21
M109 2 3 2 cpoly_p w=3.8e-06 l=2e-06 c=5.2038e-14 as=2.31158e-13 ad=7.488e-13 ps=1.44e-06 pd=1.11673e-06 sim_w=2.88e-06 m_per_maxw=1.31944 numb_sub_cont=3 nfing=1 $X=-827020 $Y=276580 $D=21
M110 2 3 2 cpoly_p w=3.8e-06 l=2e-06 c=5.2038e-14 as=2.31158e-13 ad=7.488e-13 ps=1.44e-06 pd=1.11673e-06 sim_w=2.88e-06 m_per_maxw=1.31944 numb_sub_cont=3 nfing=1 $X=-824500 $Y=276580 $D=21
M111 2 3 2 cpoly_p w=3.8e-06 l=2e-06 c=5.2038e-14 as=2.31158e-13 ad=7.488e-13 ps=1.44e-06 pd=1.11673e-06 sim_w=2.88e-06 m_per_maxw=1.31944 numb_sub_cont=3 nfing=1 $X=-821980 $Y=276580 $D=21
M112 2 3 2 cpoly_p w=3.8e-06 l=2e-06 c=5.2038e-14 as=2.31158e-13 ad=7.488e-13 ps=1.44e-06 pd=1.11673e-06 sim_w=2.88e-06 m_per_maxw=1.31944 numb_sub_cont=3 nfing=1 $X=-819460 $Y=276580 $D=21
M113 2 3 2 cpoly_p w=3.8e-06 l=2e-06 c=5.2038e-14 as=2.31158e-13 ad=7.488e-13 ps=1.44e-06 pd=1.11673e-06 sim_w=2.88e-06 m_per_maxw=1.31944 numb_sub_cont=3 nfing=1 $X=-816940 $Y=276580 $D=21
M114 2 3 2 cpoly_p w=3.8e-06 l=2e-06 c=5.2038e-14 as=2.31158e-13 ad=7.488e-13 ps=1.44e-06 pd=1.11673e-06 sim_w=2.88e-06 m_per_maxw=1.31944 numb_sub_cont=3 nfing=1 $X=-814420 $Y=276580 $D=21
M115 2 3 2 cpoly_p w=3.8e-06 l=2e-06 c=5.2038e-14 as=2.31158e-13 ad=7.488e-13 ps=1.44e-06 pd=1.11673e-06 sim_w=2.88e-06 m_per_maxw=1.31944 numb_sub_cont=3 nfing=1 $X=-811900 $Y=276580 $D=21
M116 2 3 2 cpoly_p w=3.8e-06 l=2e-06 c=5.2038e-14 as=2.31158e-13 ad=7.488e-13 ps=1.44e-06 pd=1.11673e-06 sim_w=2.88e-06 m_per_maxw=1.31944 numb_sub_cont=3 nfing=1 $X=-809380 $Y=276580 $D=21
M117 2 3 2 cpoly_p w=3.8e-06 l=2e-06 c=5.2038e-14 as=2.31158e-13 ad=7.488e-13 ps=1.44e-06 pd=1.11673e-06 sim_w=2.88e-06 m_per_maxw=1.31944 numb_sub_cont=3 nfing=1 $X=-806860 $Y=276580 $D=21
M118 2 3 2 cpoly_p w=3.8e-06 l=2e-06 c=5.2038e-14 as=2.31158e-13 ad=7.488e-13 ps=1.44e-06 pd=1.11673e-06 sim_w=2.88e-06 m_per_maxw=1.31944 numb_sub_cont=3 nfing=1 $X=-804340 $Y=276580 $D=21
M119 2 3 2 cpoly_p w=3.8e-06 l=2e-06 c=5.2038e-14 as=2.31158e-13 ad=7.488e-13 ps=1.44e-06 pd=1.11673e-06 sim_w=2.88e-06 m_per_maxw=1.31944 numb_sub_cont=3 nfing=1 $X=-801820 $Y=276580 $D=21
M120 2 3 2 cpoly_p w=3.8e-06 l=2e-06 c=5.2038e-14 as=2.31158e-13 ad=7.488e-13 ps=1.44e-06 pd=1.11673e-06 sim_w=2.88e-06 m_per_maxw=1.31944 numb_sub_cont=3 nfing=1 $X=-799300 $Y=276580 $D=21
M121 2 3 2 cpoly_p w=3.8e-06 l=2e-06 c=5.2038e-14 as=2.31158e-13 ad=7.488e-13 ps=1.44e-06 pd=1.11673e-06 sim_w=2.88e-06 m_per_maxw=1.31944 numb_sub_cont=3 nfing=1 $X=-796780 $Y=276580 $D=21
M122 2 3 2 cpoly_p w=3.8e-06 l=2e-06 c=5.2038e-14 as=2.31158e-13 ad=7.488e-13 ps=1.44e-06 pd=1.11673e-06 sim_w=2.88e-06 m_per_maxw=1.31944 numb_sub_cont=3 nfing=1 $X=-794260 $Y=276580 $D=21
M123 2 3 2 cpoly_p w=3.8e-06 l=2e-06 c=5.2038e-14 as=2.31158e-13 ad=7.488e-13 ps=1.44e-06 pd=1.11673e-06 sim_w=2.88e-06 m_per_maxw=1.31944 numb_sub_cont=3 nfing=1 $X=-791740 $Y=276580 $D=21
M124 2 3 2 cpoly_p w=3.8e-06 l=2e-06 c=5.2038e-14 as=2.31158e-13 ad=7.488e-13 ps=1.44e-06 pd=1.11673e-06 sim_w=2.88e-06 m_per_maxw=1.31944 numb_sub_cont=3 nfing=1 $X=-789220 $Y=276580 $D=21
M125 2 3 2 cpoly_p w=3.8e-06 l=2e-06 c=5.2038e-14 as=2.31158e-13 ad=7.488e-13 ps=1.44e-06 pd=1.11673e-06 sim_w=2.88e-06 m_per_maxw=1.31944 numb_sub_cont=3 nfing=1 $X=-786700 $Y=276580 $D=21
M126 2 3 2 cpoly_p w=3.8e-06 l=2e-06 c=5.2038e-14 as=2.31158e-13 ad=7.488e-13 ps=1.44e-06 pd=1.11673e-06 sim_w=2.88e-06 m_per_maxw=1.31944 numb_sub_cont=3 nfing=1 $X=-784180 $Y=276580 $D=21
M127 2 3 2 cpoly_p w=3.8e-06 l=2e-06 c=5.2038e-14 as=2.31158e-13 ad=7.488e-13 ps=1.44e-06 pd=1.11673e-06 sim_w=2.88e-06 m_per_maxw=1.31944 numb_sub_cont=3 nfing=1 $X=-781660 $Y=276580 $D=21
M128 2 3 2 cpoly_p w=3.8e-06 l=2e-06 c=5.2038e-14 as=2.31158e-13 ad=7.488e-13 ps=1.44e-06 pd=1.11673e-06 sim_w=2.88e-06 m_per_maxw=1.31944 numb_sub_cont=3 nfing=1 $X=-779140 $Y=276580 $D=21
M129 2 3 2 cpoly_p w=3.8e-06 l=2e-06 c=5.2038e-14 as=2.31158e-13 ad=7.488e-13 ps=1.44e-06 pd=1.11673e-06 sim_w=2.88e-06 m_per_maxw=1.31944 numb_sub_cont=3 nfing=1 $X=-776620 $Y=276580 $D=21
M130 2 3 2 cpoly_p w=3.8e-06 l=2e-06 c=5.2038e-14 as=2.31158e-13 ad=7.488e-13 ps=1.44e-06 pd=1.11673e-06 sim_w=2.88e-06 m_per_maxw=1.31944 numb_sub_cont=3 nfing=1 $X=-774100 $Y=276580 $D=21
M131 2 3 2 cpoly_p w=3.8e-06 l=2e-06 c=5.2038e-14 as=2.31158e-13 ad=7.488e-13 ps=1.44e-06 pd=1.11673e-06 sim_w=2.88e-06 m_per_maxw=1.31944 numb_sub_cont=3 nfing=1 $X=-771580 $Y=276580 $D=21
M132 2 3 2 cpoly_p w=3.8e-06 l=2e-06 c=5.2038e-14 as=2.31158e-13 ad=7.488e-13 ps=1.44e-06 pd=1.11673e-06 sim_w=2.88e-06 m_per_maxw=1.31944 numb_sub_cont=3 nfing=1 $X=-769060 $Y=276580 $D=21
M133 2 3 2 cpoly_p w=3.8e-06 l=2e-06 c=5.2038e-14 as=2.31158e-13 ad=7.488e-13 ps=1.44e-06 pd=1.11673e-06 sim_w=2.88e-06 m_per_maxw=1.31944 numb_sub_cont=3 nfing=1 $X=-766540 $Y=276580 $D=21
M134 2 3 2 cpoly_p w=3.8e-06 l=2e-06 c=5.2038e-14 as=2.31158e-13 ad=7.488e-13 ps=1.44e-06 pd=1.11673e-06 sim_w=2.88e-06 m_per_maxw=1.31944 numb_sub_cont=3 nfing=1 $X=-764020 $Y=276580 $D=21
M135 2 3 2 cpoly_p w=3.8e-06 l=2e-06 c=5.2038e-14 as=2.31158e-13 ad=7.488e-13 ps=1.44e-06 pd=1.11673e-06 sim_w=2.88e-06 m_per_maxw=1.31944 numb_sub_cont=3 nfing=1 $X=-761500 $Y=276580 $D=21
M136 2 3 2 cpoly_p w=3.8e-06 l=2e-06 c=5.2038e-14 as=2.31158e-13 ad=7.488e-13 ps=1.44e-06 pd=1.11673e-06 sim_w=2.88e-06 m_per_maxw=1.31944 numb_sub_cont=3 nfing=1 $X=-758980 $Y=276580 $D=21
M137 2 3 2 cpoly_p w=3.8e-06 l=2e-06 c=5.2038e-14 as=2.31158e-13 ad=7.488e-13 ps=1.44e-06 pd=1.11673e-06 sim_w=2.88e-06 m_per_maxw=1.31944 numb_sub_cont=3 nfing=1 $X=-756460 $Y=276580 $D=21
M138 2 3 2 cpoly_p w=3.8e-06 l=2e-06 c=5.2038e-14 as=2.31158e-13 ad=7.488e-13 ps=1.44e-06 pd=1.11673e-06 sim_w=2.88e-06 m_per_maxw=1.31944 numb_sub_cont=3 nfing=1 $X=-753940 $Y=276580 $D=21
M139 2 3 2 cpoly_p w=3.8e-06 l=2e-06 c=5.2038e-14 as=2.31158e-13 ad=7.488e-13 ps=1.44e-06 pd=1.11673e-06 sim_w=2.88e-06 m_per_maxw=1.31944 numb_sub_cont=3 nfing=1 $X=-751420 $Y=276580 $D=21
M140 2 3 2 cpoly_p w=3.8e-06 l=2e-06 c=5.2038e-14 as=2.31158e-13 ad=7.488e-13 ps=1.44e-06 pd=1.11673e-06 sim_w=2.88e-06 m_per_maxw=1.31944 numb_sub_cont=3 nfing=1 $X=-748900 $Y=276580 $D=21
M141 2 3 2 cpoly_p w=3.8e-06 l=2e-06 c=5.2038e-14 as=2.31158e-13 ad=7.488e-13 ps=1.44e-06 pd=1.11673e-06 sim_w=2.88e-06 m_per_maxw=1.31944 numb_sub_cont=3 nfing=1 $X=-746380 $Y=276580 $D=21
M142 2 3 2 cpoly_p w=3.8e-06 l=2e-06 c=5.2038e-14 as=2.31158e-13 ad=7.488e-13 ps=1.44e-06 pd=1.11673e-06 sim_w=2.88e-06 m_per_maxw=1.31944 numb_sub_cont=3 nfing=1 $X=-743860 $Y=276580 $D=21
M143 2 3 2 cpoly_p w=3.8e-06 l=2e-06 c=5.2038e-14 as=2.31158e-13 ad=7.488e-13 ps=1.44e-06 pd=1.11673e-06 sim_w=2.88e-06 m_per_maxw=1.31944 numb_sub_cont=3 nfing=1 $X=-741340 $Y=276580 $D=21
M144 2 3 2 cpoly_p w=3.8e-06 l=2e-06 c=5.2038e-14 as=2.31158e-13 ad=7.488e-13 ps=1.44e-06 pd=1.11673e-06 sim_w=2.88e-06 m_per_maxw=1.31944 numb_sub_cont=3 nfing=1 $X=-738820 $Y=276580 $D=21
M145 2 3 2 cpoly_p w=3.8e-06 l=2e-06 c=5.2038e-14 as=2.31158e-13 ad=7.488e-13 ps=1.44e-06 pd=1.11673e-06 sim_w=2.88e-06 m_per_maxw=1.31944 numb_sub_cont=3 nfing=1 $X=-736300 $Y=276580 $D=21
M146 2 3 2 cpoly_p w=3.8e-06 l=2e-06 c=5.2038e-14 as=2.31158e-13 ad=7.488e-13 ps=1.44e-06 pd=1.11673e-06 sim_w=2.88e-06 m_per_maxw=1.31944 numb_sub_cont=3 nfing=1 $X=-733780 $Y=276580 $D=21
M147 2 3 2 cpoly_p w=3.8e-06 l=2e-06 c=5.2038e-14 as=2.31158e-13 ad=7.488e-13 ps=1.44e-06 pd=1.11673e-06 sim_w=2.88e-06 m_per_maxw=1.31944 numb_sub_cont=3 nfing=1 $X=-731260 $Y=276580 $D=21
M148 2 3 2 cpoly_p w=3.8e-06 l=2e-06 c=5.2038e-14 as=2.31158e-13 ad=7.488e-13 ps=1.44e-06 pd=1.11673e-06 sim_w=2.88e-06 m_per_maxw=1.31944 numb_sub_cont=3 nfing=1 $X=-728740 $Y=276580 $D=21
M149 2 3 2 cpoly_p w=3.8e-06 l=2e-06 c=5.2038e-14 as=2.31158e-13 ad=7.488e-13 ps=1.44e-06 pd=1.11673e-06 sim_w=2.88e-06 m_per_maxw=1.31944 numb_sub_cont=3 nfing=1 $X=-726220 $Y=276580 $D=21
M150 2 3 2 cpoly_p w=3.8e-06 l=2e-06 c=5.2038e-14 as=2.31158e-13 ad=7.488e-13 ps=1.44e-06 pd=1.11673e-06 sim_w=2.88e-06 m_per_maxw=1.31944 numb_sub_cont=3 nfing=1 $X=-723700 $Y=276580 $D=21
M151 2 3 2 cpoly_p w=3.8e-06 l=2e-06 c=5.2038e-14 as=2.31158e-13 ad=7.488e-13 ps=1.44e-06 pd=1.11673e-06 sim_w=2.88e-06 m_per_maxw=1.31944 numb_sub_cont=3 nfing=1 $X=-721180 $Y=276580 $D=21
M152 2 3 2 cpoly_p w=3.8e-06 l=2e-06 c=5.2038e-14 as=2.31158e-13 ad=7.488e-13 ps=1.44e-06 pd=1.11673e-06 sim_w=2.88e-06 m_per_maxw=1.31944 numb_sub_cont=3 nfing=1 $X=-718660 $Y=276580 $D=21
M153 2 3 2 cpoly_p w=3.8e-06 l=2e-06 c=5.2038e-14 as=2.31158e-13 ad=7.488e-13 ps=1.44e-06 pd=1.11673e-06 sim_w=2.88e-06 m_per_maxw=1.31944 numb_sub_cont=3 nfing=1 $X=-716140 $Y=276580 $D=21
M154 2 3 2 cpoly_p w=3.8e-06 l=2e-06 c=5.2038e-14 as=2.31158e-13 ad=7.488e-13 ps=1.44e-06 pd=1.11673e-06 sim_w=2.88e-06 m_per_maxw=1.31944 numb_sub_cont=3 nfing=1 $X=-713620 $Y=276580 $D=21
M155 2 3 2 cpoly_p w=3.8e-06 l=2e-06 c=5.2038e-14 as=2.31158e-13 ad=7.488e-13 ps=1.44e-06 pd=1.11673e-06 sim_w=2.88e-06 m_per_maxw=1.31944 numb_sub_cont=3 nfing=1 $X=-711100 $Y=276580 $D=21
M156 2 3 2 cpoly_p w=3.8e-06 l=2e-06 c=5.2038e-14 as=2.31158e-13 ad=7.488e-13 ps=1.44e-06 pd=1.11673e-06 sim_w=2.88e-06 m_per_maxw=1.31944 numb_sub_cont=3 nfing=1 $X=-708580 $Y=276580 $D=21
M157 2 3 2 cpoly_p w=3.8e-06 l=2e-06 c=5.2038e-14 as=2.31158e-13 ad=7.488e-13 ps=1.44e-06 pd=1.11673e-06 sim_w=2.88e-06 m_per_maxw=1.31944 numb_sub_cont=3 nfing=1 $X=-706060 $Y=276580 $D=21
M158 2 3 2 cpoly_p w=3.8e-06 l=2e-06 c=5.2038e-14 as=2.31158e-13 ad=7.488e-13 ps=1.44e-06 pd=1.11673e-06 sim_w=2.88e-06 m_per_maxw=1.31944 numb_sub_cont=3 nfing=1 $X=-703540 $Y=276580 $D=21
M159 2 3 2 cpoly_p w=3.8e-06 l=2e-06 c=5.2038e-14 as=2.31158e-13 ad=7.488e-13 ps=1.44e-06 pd=1.11673e-06 sim_w=2.88e-06 m_per_maxw=1.31944 numb_sub_cont=3 nfing=1 $X=-701020 $Y=276580 $D=21
M160 2 3 2 cpoly_p w=3.8e-06 l=2e-06 c=5.2038e-14 as=2.31158e-13 ad=7.488e-13 ps=1.44e-06 pd=1.11673e-06 sim_w=2.88e-06 m_per_maxw=1.31944 numb_sub_cont=3 nfing=1 $X=-698500 $Y=276580 $D=21
M161 2 3 2 cpoly_p w=3.8e-06 l=2e-06 c=5.2038e-14 as=2.31158e-13 ad=7.488e-13 ps=1.44e-06 pd=1.11673e-06 sim_w=2.88e-06 m_per_maxw=1.31944 numb_sub_cont=3 nfing=1 $X=-695980 $Y=276580 $D=21
M162 2 3 2 cpoly_p w=3.8e-06 l=2e-06 c=5.2038e-14 as=2.31158e-13 ad=7.488e-13 ps=1.44e-06 pd=1.11673e-06 sim_w=2.88e-06 m_per_maxw=1.31944 numb_sub_cont=3 nfing=1 $X=-693460 $Y=276580 $D=21
M163 2 3 2 cpoly_p w=3.8e-06 l=2e-06 c=5.2038e-14 as=2.31158e-13 ad=7.488e-13 ps=1.44e-06 pd=1.11673e-06 sim_w=2.88e-06 m_per_maxw=1.31944 numb_sub_cont=3 nfing=1 $X=-690940 $Y=276580 $D=21
M164 2 3 2 cpoly_p w=3.8e-06 l=2e-06 c=5.2038e-14 as=2.31158e-13 ad=7.488e-13 ps=1.44e-06 pd=1.11673e-06 sim_w=2.88e-06 m_per_maxw=1.31944 numb_sub_cont=3 nfing=1 $X=-688420 $Y=276580 $D=21
M165 2 3 2 cpoly_p w=3.8e-06 l=2e-06 c=5.2038e-14 as=2.31158e-13 ad=7.488e-13 ps=1.44e-06 pd=1.11673e-06 sim_w=2.88e-06 m_per_maxw=1.31944 numb_sub_cont=3 nfing=1 $X=-685900 $Y=276580 $D=21
M166 2 3 2 cpoly_p w=3.8e-06 l=2e-06 c=5.2038e-14 as=2.31158e-13 ad=7.488e-13 ps=1.44e-06 pd=1.11673e-06 sim_w=2.88e-06 m_per_maxw=1.31944 numb_sub_cont=3 nfing=1 $X=-683380 $Y=276580 $D=21
M167 2 3 2 cpoly_p w=3.8e-06 l=2e-06 c=5.2038e-14 as=2.31158e-13 ad=7.488e-13 ps=1.44e-06 pd=1.11673e-06 sim_w=2.88e-06 m_per_maxw=1.31944 numb_sub_cont=3 nfing=1 $X=-680860 $Y=276580 $D=21
M168 2 3 2 cpoly_p w=3.8e-06 l=2e-06 c=5.2038e-14 as=2.31158e-13 ad=7.488e-13 ps=1.44e-06 pd=1.11673e-06 sim_w=2.88e-06 m_per_maxw=1.31944 numb_sub_cont=3 nfing=1 $X=-678340 $Y=276580 $D=21
M169 2 3 2 cpoly_p w=3.8e-06 l=2e-06 c=5.2038e-14 as=2.31158e-13 ad=7.488e-13 ps=1.44e-06 pd=1.11673e-06 sim_w=2.88e-06 m_per_maxw=1.31944 numb_sub_cont=3 nfing=1 $X=-675820 $Y=276580 $D=21
M170 2 3 2 cpoly_p w=3.8e-06 l=2e-06 c=5.2038e-14 as=2.31158e-13 ad=7.488e-13 ps=1.44e-06 pd=1.11673e-06 sim_w=2.88e-06 m_per_maxw=1.31944 numb_sub_cont=3 nfing=1 $X=-673300 $Y=276580 $D=21
M171 2 3 2 cpoly_p w=3.8e-06 l=2e-06 c=5.2038e-14 as=2.31158e-13 ad=7.488e-13 ps=1.44e-06 pd=1.11673e-06 sim_w=2.88e-06 m_per_maxw=1.31944 numb_sub_cont=3 nfing=1 $X=-670780 $Y=276580 $D=21
M172 2 3 2 cpoly_p w=3.8e-06 l=2e-06 c=5.2038e-14 as=2.31158e-13 ad=7.488e-13 ps=1.44e-06 pd=1.11673e-06 sim_w=2.88e-06 m_per_maxw=1.31944 numb_sub_cont=3 nfing=1 $X=-668260 $Y=276580 $D=21
M173 2 3 2 cpoly_p w=3.8e-06 l=2e-06 c=5.2038e-14 as=2.31158e-13 ad=7.488e-13 ps=1.44e-06 pd=1.11673e-06 sim_w=2.88e-06 m_per_maxw=1.31944 numb_sub_cont=3 nfing=1 $X=-665740 $Y=276580 $D=21
M174 2 3 2 cpoly_p w=3.8e-06 l=2e-06 c=5.2038e-14 as=2.31158e-13 ad=7.488e-13 ps=1.44e-06 pd=1.11673e-06 sim_w=2.88e-06 m_per_maxw=1.31944 numb_sub_cont=3 nfing=1 $X=-663220 $Y=276580 $D=21
M175 2 3 2 cpoly_p w=3.8e-06 l=2e-06 c=5.2038e-14 as=2.31158e-13 ad=7.488e-13 ps=1.44e-06 pd=1.11673e-06 sim_w=2.88e-06 m_per_maxw=1.31944 numb_sub_cont=3 nfing=1 $X=-660700 $Y=276580 $D=21
M176 2 3 2 cpoly_p w=3.8e-06 l=2e-06 c=5.2038e-14 as=2.31158e-13 ad=7.488e-13 ps=1.44e-06 pd=1.11673e-06 sim_w=2.88e-06 m_per_maxw=1.31944 numb_sub_cont=3 nfing=1 $X=-658180 $Y=276580 $D=21
M177 2 3 2 cpoly_p w=3.8e-06 l=2e-06 c=5.2038e-14 as=2.31158e-13 ad=7.488e-13 ps=1.44e-06 pd=1.11673e-06 sim_w=2.88e-06 m_per_maxw=1.31944 numb_sub_cont=3 nfing=1 $X=-655660 $Y=276580 $D=21
M178 2 3 2 cpoly_p w=3.8e-06 l=2e-06 c=5.2038e-14 as=2.31158e-13 ad=7.488e-13 ps=1.44e-06 pd=1.11673e-06 sim_w=2.88e-06 m_per_maxw=1.31944 numb_sub_cont=3 nfing=1 $X=-653140 $Y=276580 $D=21
M179 2 3 2 cpoly_p w=3.8e-06 l=2e-06 c=5.2038e-14 as=2.31158e-13 ad=7.488e-13 ps=1.44e-06 pd=1.11673e-06 sim_w=2.88e-06 m_per_maxw=1.31944 numb_sub_cont=3 nfing=1 $X=-650620 $Y=276580 $D=21
M180 2 3 2 cpoly_p w=3.8e-06 l=2e-06 c=5.2038e-14 as=2.31158e-13 ad=7.488e-13 ps=1.44e-06 pd=1.11673e-06 sim_w=2.88e-06 m_per_maxw=1.31944 numb_sub_cont=3 nfing=1 $X=-648100 $Y=276580 $D=21
M181 2 3 2 cpoly_p w=3.8e-06 l=2e-06 c=5.2038e-14 as=2.31158e-13 ad=7.488e-13 ps=1.44e-06 pd=1.11673e-06 sim_w=2.88e-06 m_per_maxw=1.31944 numb_sub_cont=3 nfing=1 $X=-645580 $Y=276580 $D=21
M182 2 3 2 cpoly_p w=3.8e-06 l=2e-06 c=5.2038e-14 as=2.31158e-13 ad=7.488e-13 ps=1.44e-06 pd=1.11673e-06 sim_w=2.88e-06 m_per_maxw=1.31944 numb_sub_cont=3 nfing=1 $X=-643060 $Y=276580 $D=21
M183 2 3 2 cpoly_p w=3.8e-06 l=2e-06 c=5.2038e-14 as=2.31158e-13 ad=7.488e-13 ps=1.44e-06 pd=1.11673e-06 sim_w=2.88e-06 m_per_maxw=1.31944 numb_sub_cont=3 nfing=1 $X=-640540 $Y=276580 $D=21
M184 2 3 2 cpoly_p w=3.8e-06 l=2e-06 c=5.2038e-14 as=2.31158e-13 ad=7.488e-13 ps=1.44e-06 pd=1.11673e-06 sim_w=2.88e-06 m_per_maxw=1.31944 numb_sub_cont=3 nfing=1 $X=-638020 $Y=276580 $D=21
M185 2 3 2 cpoly_p w=3.8e-06 l=2e-06 c=5.2038e-14 as=2.31158e-13 ad=7.488e-13 ps=1.44e-06 pd=1.11673e-06 sim_w=2.88e-06 m_per_maxw=1.31944 numb_sub_cont=3 nfing=1 $X=-635500 $Y=276580 $D=21
M186 2 3 2 cpoly_p w=3.8e-06 l=2e-06 c=5.2038e-14 as=2.31158e-13 ad=7.488e-13 ps=1.44e-06 pd=1.11673e-06 sim_w=2.88e-06 m_per_maxw=1.31944 numb_sub_cont=3 nfing=1 $X=-632980 $Y=276580 $D=21
M187 2 3 2 cpoly_p w=3.8e-06 l=2e-06 c=5.2038e-14 as=2.31158e-13 ad=7.488e-13 ps=1.44e-06 pd=1.11673e-06 sim_w=2.88e-06 m_per_maxw=1.31944 numb_sub_cont=3 nfing=1 $X=-630460 $Y=276580 $D=21
M188 2 3 2 cpoly_p w=3.8e-06 l=2e-06 c=5.2038e-14 as=2.31158e-13 ad=7.488e-13 ps=1.44e-06 pd=1.11673e-06 sim_w=2.88e-06 m_per_maxw=1.31944 numb_sub_cont=3 nfing=1 $X=-627940 $Y=276580 $D=21
M189 2 3 2 cpoly_p w=3.8e-06 l=2e-06 c=5.2038e-14 as=2.31158e-13 ad=7.488e-13 ps=1.44e-06 pd=1.11673e-06 sim_w=2.88e-06 m_per_maxw=1.31944 numb_sub_cont=3 nfing=1 $X=-625420 $Y=276580 $D=21
M190 2 3 2 cpoly_p w=3.8e-06 l=2e-06 c=5.2038e-14 as=2.31158e-13 ad=7.488e-13 ps=1.44e-06 pd=1.11673e-06 sim_w=2.88e-06 m_per_maxw=1.31944 numb_sub_cont=3 nfing=1 $X=-622900 $Y=276580 $D=21
M191 2 3 2 cpoly_p w=3.8e-06 l=2e-06 c=5.2038e-14 as=2.31158e-13 ad=7.488e-13 ps=1.44e-06 pd=1.11673e-06 sim_w=2.88e-06 m_per_maxw=1.31944 numb_sub_cont=3 nfing=1 $X=-620380 $Y=276580 $D=21
M192 2 3 2 cpoly_p w=3.8e-06 l=2e-06 c=5.2038e-14 as=2.31158e-13 ad=7.488e-13 ps=1.44e-06 pd=1.11673e-06 sim_w=2.88e-06 m_per_maxw=1.31944 numb_sub_cont=3 nfing=1 $X=-617860 $Y=276580 $D=21
M193 2 3 2 cpoly_p w=3.8e-06 l=2e-06 c=5.2038e-14 as=2.31158e-13 ad=7.488e-13 ps=1.44e-06 pd=1.11673e-06 sim_w=2.88e-06 m_per_maxw=1.31944 numb_sub_cont=3 nfing=1 $X=-615340 $Y=276580 $D=21
M194 2 3 2 cpoly_p w=3.8e-06 l=2e-06 c=5.2038e-14 as=2.31158e-13 ad=7.488e-13 ps=1.44e-06 pd=1.11673e-06 sim_w=2.88e-06 m_per_maxw=1.31944 numb_sub_cont=3 nfing=1 $X=-612820 $Y=276580 $D=21
M195 2 3 2 cpoly_p w=3.8e-06 l=2e-06 c=5.2038e-14 as=2.31158e-13 ad=7.488e-13 ps=1.44e-06 pd=1.11673e-06 sim_w=2.88e-06 m_per_maxw=1.31944 numb_sub_cont=3 nfing=1 $X=-610300 $Y=276580 $D=21
M196 2 3 2 cpoly_p w=3.8e-06 l=2e-06 c=5.2038e-14 as=2.31158e-13 ad=7.488e-13 ps=1.44e-06 pd=1.11673e-06 sim_w=2.88e-06 m_per_maxw=1.31944 numb_sub_cont=3 nfing=1 $X=-607780 $Y=276580 $D=21
M197 2 3 2 cpoly_p w=3.8e-06 l=2e-06 c=5.2038e-14 as=2.31158e-13 ad=7.488e-13 ps=1.44e-06 pd=1.11673e-06 sim_w=2.88e-06 m_per_maxw=1.31944 numb_sub_cont=3 nfing=1 $X=-605260 $Y=276580 $D=21
M198 2 3 2 cpoly_p w=3.8e-06 l=2e-06 c=5.2038e-14 as=2.31158e-13 ad=7.488e-13 ps=1.44e-06 pd=1.11673e-06 sim_w=2.88e-06 m_per_maxw=1.31944 numb_sub_cont=3 nfing=1 $X=-602740 $Y=276580 $D=21
M199 2 3 2 cpoly_p w=3.8e-06 l=2e-06 c=5.2038e-14 as=2.31158e-13 ad=7.488e-13 ps=1.44e-06 pd=1.11673e-06 sim_w=2.88e-06 m_per_maxw=1.31944 numb_sub_cont=3 nfing=1 $X=-600220 $Y=276580 $D=21
M200 2 3 2 cpoly_p w=3.8e-06 l=2e-06 c=5.2038e-14 as=2.31158e-13 ad=7.488e-13 ps=1.44e-06 pd=1.11673e-06 sim_w=2.88e-06 m_per_maxw=1.31944 numb_sub_cont=3 nfing=1 $X=-597700 $Y=276580 $D=21
M201 2 3 2 cpoly_p w=3.8e-06 l=2e-06 c=5.2038e-14 as=2.31158e-13 ad=7.488e-13 ps=1.44e-06 pd=1.11673e-06 sim_w=2.88e-06 m_per_maxw=1.31944 numb_sub_cont=3 nfing=1 $X=-595180 $Y=276580 $D=21
M202 2 3 2 cpoly_p w=3.8e-06 l=2e-06 c=5.2038e-14 as=2.31158e-13 ad=7.488e-13 ps=1.44e-06 pd=1.11673e-06 sim_w=2.88e-06 m_per_maxw=1.31944 numb_sub_cont=3 nfing=1 $X=-592660 $Y=276580 $D=21
M203 2 3 2 cpoly_p w=3.8e-06 l=2e-06 c=5.2038e-14 as=2.31158e-13 ad=7.488e-13 ps=1.44e-06 pd=1.11673e-06 sim_w=2.88e-06 m_per_maxw=1.31944 numb_sub_cont=3 nfing=1 $X=-590140 $Y=276580 $D=21
M204 2 3 2 cpoly_p w=3.8e-06 l=2e-06 c=5.2038e-14 as=2.31158e-13 ad=7.488e-13 ps=1.44e-06 pd=1.11673e-06 sim_w=2.88e-06 m_per_maxw=1.31944 numb_sub_cont=3 nfing=1 $X=-587620 $Y=276580 $D=21
M205 2 3 2 cpoly_p w=3.8e-06 l=2e-06 c=5.2038e-14 as=2.31158e-13 ad=7.488e-13 ps=1.44e-06 pd=1.11673e-06 sim_w=2.88e-06 m_per_maxw=1.31944 numb_sub_cont=3 nfing=1 $X=-585100 $Y=276580 $D=21
M206 2 3 2 cpoly_p w=3.8e-06 l=2e-06 c=5.2038e-14 as=2.31158e-13 ad=7.488e-13 ps=1.44e-06 pd=1.11673e-06 sim_w=2.88e-06 m_per_maxw=1.31944 numb_sub_cont=3 nfing=1 $X=-582580 $Y=276580 $D=21
M207 2 3 2 cpoly_p w=3.8e-06 l=2e-06 c=5.2038e-14 as=2.31158e-13 ad=7.488e-13 ps=1.44e-06 pd=1.11673e-06 sim_w=2.88e-06 m_per_maxw=1.31944 numb_sub_cont=3 nfing=1 $X=-580060 $Y=276580 $D=21
M208 2 3 2 cpoly_p w=3.8e-06 l=2e-06 c=5.2038e-14 as=2.31158e-13 ad=7.488e-13 ps=1.44e-06 pd=1.11673e-06 sim_w=2.88e-06 m_per_maxw=1.31944 numb_sub_cont=3 nfing=1 $X=-577540 $Y=276580 $D=21
M209 2 3 2 cpoly_p w=3.8e-06 l=2e-06 c=5.2038e-14 as=2.31158e-13 ad=7.488e-13 ps=1.44e-06 pd=1.11673e-06 sim_w=2.88e-06 m_per_maxw=1.31944 numb_sub_cont=3 nfing=1 $X=-575020 $Y=276580 $D=21
M210 2 3 2 cpoly_p w=3.8e-06 l=2e-06 c=5.2038e-14 as=2.31158e-13 ad=7.488e-13 ps=1.44e-06 pd=1.11673e-06 sim_w=2.88e-06 m_per_maxw=1.31944 numb_sub_cont=3 nfing=1 $X=-572500 $Y=276580 $D=21
M211 2 3 2 cpoly_p w=3.8e-06 l=2e-06 c=5.2038e-14 as=2.31158e-13 ad=7.488e-13 ps=1.44e-06 pd=1.11673e-06 sim_w=2.88e-06 m_per_maxw=1.31944 numb_sub_cont=3 nfing=1 $X=-569980 $Y=276580 $D=21
M212 2 3 2 cpoly_p w=3.8e-06 l=2e-06 c=5.2038e-14 as=2.31158e-13 ad=7.488e-13 ps=1.44e-06 pd=1.11673e-06 sim_w=2.88e-06 m_per_maxw=1.31944 numb_sub_cont=3 nfing=1 $X=-567460 $Y=276580 $D=21
M213 2 3 2 cpoly_p w=3.8e-06 l=2e-06 c=5.2038e-14 as=2.31158e-13 ad=7.488e-13 ps=1.44e-06 pd=1.11673e-06 sim_w=2.88e-06 m_per_maxw=1.31944 numb_sub_cont=3 nfing=1 $X=-564940 $Y=276580 $D=21
M214 2 3 2 cpoly_p w=3.8e-06 l=2e-06 c=5.2038e-14 as=2.31158e-13 ad=7.488e-13 ps=1.44e-06 pd=1.11673e-06 sim_w=2.88e-06 m_per_maxw=1.31944 numb_sub_cont=3 nfing=1 $X=-562420 $Y=276580 $D=21
M215 2 3 2 cpoly_p w=3.8e-06 l=2e-06 c=5.2038e-14 as=2.31158e-13 ad=7.488e-13 ps=1.44e-06 pd=1.11673e-06 sim_w=2.88e-06 m_per_maxw=1.31944 numb_sub_cont=3 nfing=1 $X=-559900 $Y=276580 $D=21
M216 2 3 2 cpoly_p w=3.8e-06 l=2e-06 c=5.2038e-14 as=2.31158e-13 ad=7.488e-13 ps=1.44e-06 pd=1.11673e-06 sim_w=2.88e-06 m_per_maxw=1.31944 numb_sub_cont=3 nfing=1 $X=-557380 $Y=276580 $D=21
M217 2 3 2 cpoly_p w=3.8e-06 l=2e-06 c=5.2038e-14 as=2.31158e-13 ad=7.488e-13 ps=1.44e-06 pd=1.11673e-06 sim_w=2.88e-06 m_per_maxw=1.31944 numb_sub_cont=3 nfing=1 $X=-554860 $Y=276580 $D=21
M218 2 3 2 cpoly_p w=3.8e-06 l=2e-06 c=5.2038e-14 as=2.31158e-13 ad=7.488e-13 ps=1.44e-06 pd=1.11673e-06 sim_w=2.88e-06 m_per_maxw=1.31944 numb_sub_cont=3 nfing=1 $X=-552340 $Y=276580 $D=21
M219 2 3 2 cpoly_p w=3.8e-06 l=2e-06 c=5.2038e-14 as=2.31158e-13 ad=7.488e-13 ps=1.44e-06 pd=1.11673e-06 sim_w=2.88e-06 m_per_maxw=1.31944 numb_sub_cont=3 nfing=1 $X=-549820 $Y=276580 $D=21
M220 2 3 2 cpoly_p w=3.8e-06 l=2e-06 c=5.2038e-14 as=2.31158e-13 ad=7.488e-13 ps=1.44e-06 pd=1.11673e-06 sim_w=2.88e-06 m_per_maxw=1.31944 numb_sub_cont=3 nfing=1 $X=-547300 $Y=276580 $D=21
M221 2 3 2 cpoly_p w=3.8e-06 l=2e-06 c=5.2038e-14 as=2.31158e-13 ad=7.488e-13 ps=1.44e-06 pd=1.11673e-06 sim_w=2.88e-06 m_per_maxw=1.31944 numb_sub_cont=3 nfing=1 $X=-544780 $Y=276580 $D=21
M222 2 3 2 cpoly_p w=3.8e-06 l=2e-06 c=5.2038e-14 as=2.31158e-13 ad=7.488e-13 ps=1.44e-06 pd=1.11673e-06 sim_w=2.88e-06 m_per_maxw=1.31944 numb_sub_cont=3 nfing=1 $X=-542260 $Y=276580 $D=21
M223 2 3 2 cpoly_p w=3.8e-06 l=2e-06 c=5.2038e-14 as=2.31158e-13 ad=7.488e-13 ps=1.44e-06 pd=1.11673e-06 sim_w=2.88e-06 m_per_maxw=1.31944 numb_sub_cont=3 nfing=1 $X=-539740 $Y=276580 $D=21
M224 2 3 2 cpoly_p w=3.8e-06 l=2e-06 c=5.2038e-14 as=2.31158e-13 ad=7.488e-13 ps=1.44e-06 pd=1.11673e-06 sim_w=2.88e-06 m_per_maxw=1.31944 numb_sub_cont=3 nfing=1 $X=-537220 $Y=276580 $D=21
M225 2 3 2 cpoly_p w=3.8e-06 l=2e-06 c=5.2038e-14 as=2.31158e-13 ad=7.488e-13 ps=1.44e-06 pd=1.11673e-06 sim_w=2.88e-06 m_per_maxw=1.31944 numb_sub_cont=3 nfing=1 $X=-534700 $Y=276580 $D=21
M226 2 3 2 cpoly_p w=3.8e-06 l=2e-06 c=5.2038e-14 as=2.31158e-13 ad=7.488e-13 ps=1.44e-06 pd=1.11673e-06 sim_w=2.88e-06 m_per_maxw=1.31944 numb_sub_cont=3 nfing=1 $X=-532180 $Y=276580 $D=21
M227 2 3 2 cpoly_p w=3.8e-06 l=2e-06 c=5.2038e-14 as=2.31158e-13 ad=7.488e-13 ps=1.44e-06 pd=1.11673e-06 sim_w=2.88e-06 m_per_maxw=1.31944 numb_sub_cont=3 nfing=1 $X=-529660 $Y=276580 $D=21
M228 2 3 2 cpoly_p w=3.8e-06 l=2e-06 c=5.2038e-14 as=2.31158e-13 ad=7.488e-13 ps=1.44e-06 pd=1.11673e-06 sim_w=2.88e-06 m_per_maxw=1.31944 numb_sub_cont=3 nfing=1 $X=-527140 $Y=276580 $D=21
M229 2 3 2 cpoly_p w=3.8e-06 l=2e-06 c=5.2038e-14 as=2.31158e-13 ad=7.488e-13 ps=1.44e-06 pd=1.11673e-06 sim_w=2.88e-06 m_per_maxw=1.31944 numb_sub_cont=3 nfing=1 $X=-524620 $Y=276580 $D=21
M230 2 3 2 cpoly_p w=3.8e-06 l=2e-06 c=5.2038e-14 as=2.31158e-13 ad=7.488e-13 ps=1.44e-06 pd=1.11673e-06 sim_w=2.88e-06 m_per_maxw=1.31944 numb_sub_cont=3 nfing=1 $X=-522100 $Y=276580 $D=21
M231 2 3 2 cpoly_p w=3.8e-06 l=2e-06 c=5.2038e-14 as=2.31158e-13 ad=7.488e-13 ps=1.44e-06 pd=1.11673e-06 sim_w=2.88e-06 m_per_maxw=1.31944 numb_sub_cont=3 nfing=1 $X=-519580 $Y=276580 $D=21
M232 2 3 2 cpoly_p w=3.8e-06 l=2e-06 c=5.2038e-14 as=2.31158e-13 ad=7.488e-13 ps=1.44e-06 pd=1.11673e-06 sim_w=2.88e-06 m_per_maxw=1.31944 numb_sub_cont=3 nfing=1 $X=-517060 $Y=276580 $D=21
M233 2 3 2 cpoly_p w=3.8e-06 l=2e-06 c=5.2038e-14 as=2.31158e-13 ad=7.488e-13 ps=1.44e-06 pd=1.11673e-06 sim_w=2.88e-06 m_per_maxw=1.31944 numb_sub_cont=3 nfing=1 $X=-514540 $Y=276580 $D=21
M234 2 3 2 cpoly_p w=3.8e-06 l=2e-06 c=5.2038e-14 as=2.31158e-13 ad=7.488e-13 ps=1.44e-06 pd=1.11673e-06 sim_w=2.88e-06 m_per_maxw=1.31944 numb_sub_cont=3 nfing=1 $X=-512020 $Y=276580 $D=21
M235 2 3 2 cpoly_p w=3.8e-06 l=2e-06 c=5.2038e-14 as=2.31158e-13 ad=7.488e-13 ps=1.44e-06 pd=1.11673e-06 sim_w=2.88e-06 m_per_maxw=1.31944 numb_sub_cont=3 nfing=1 $X=-509500 $Y=276580 $D=21
M236 2 3 2 cpoly_p w=3.8e-06 l=2e-06 c=5.2038e-14 as=2.31158e-13 ad=7.488e-13 ps=1.44e-06 pd=1.11673e-06 sim_w=2.88e-06 m_per_maxw=1.31944 numb_sub_cont=3 nfing=1 $X=-506980 $Y=276580 $D=21
M237 2 3 2 cpoly_p w=3.8e-06 l=2e-06 c=5.2038e-14 as=2.31158e-13 ad=7.488e-13 ps=1.44e-06 pd=1.11673e-06 sim_w=2.88e-06 m_per_maxw=1.31944 numb_sub_cont=3 nfing=1 $X=-504460 $Y=276580 $D=21
M238 2 3 2 cpoly_p w=3.8e-06 l=2e-06 c=5.2038e-14 as=2.31158e-13 ad=7.488e-13 ps=1.44e-06 pd=1.11673e-06 sim_w=2.88e-06 m_per_maxw=1.31944 numb_sub_cont=3 nfing=1 $X=-501940 $Y=276580 $D=21
M239 2 3 2 cpoly_p w=3.8e-06 l=2e-06 c=5.2038e-14 as=2.31158e-13 ad=7.488e-13 ps=1.44e-06 pd=1.11673e-06 sim_w=2.88e-06 m_per_maxw=1.31944 numb_sub_cont=3 nfing=1 $X=-499420 $Y=276580 $D=21
M240 2 3 2 cpoly_p w=3.8e-06 l=2e-06 c=5.2038e-14 as=2.31158e-13 ad=7.488e-13 ps=1.44e-06 pd=1.11673e-06 sim_w=2.88e-06 m_per_maxw=1.31944 numb_sub_cont=3 nfing=1 $X=-496900 $Y=276580 $D=21
M241 2 3 2 cpoly_p w=3.8e-06 l=2e-06 c=5.2038e-14 as=2.31158e-13 ad=7.488e-13 ps=1.44e-06 pd=1.11673e-06 sim_w=2.88e-06 m_per_maxw=1.31944 numb_sub_cont=3 nfing=1 $X=-494380 $Y=276580 $D=21
M242 2 3 2 cpoly_p w=3.8e-06 l=2e-06 c=5.2038e-14 as=2.31158e-13 ad=7.488e-13 ps=1.44e-06 pd=1.11673e-06 sim_w=2.88e-06 m_per_maxw=1.31944 numb_sub_cont=3 nfing=1 $X=-491860 $Y=276580 $D=21
M243 2 3 2 cpoly_p w=3.8e-06 l=2e-06 c=5.2038e-14 as=2.31158e-13 ad=7.488e-13 ps=1.44e-06 pd=1.11673e-06 sim_w=2.88e-06 m_per_maxw=1.31944 numb_sub_cont=3 nfing=1 $X=-489340 $Y=276580 $D=21
M244 2 3 2 cpoly_p w=3.8e-06 l=2e-06 c=5.2038e-14 as=2.31158e-13 ad=7.488e-13 ps=1.44e-06 pd=1.11673e-06 sim_w=2.88e-06 m_per_maxw=1.31944 numb_sub_cont=3 nfing=1 $X=-486820 $Y=276580 $D=21
M245 2 3 2 cpoly_p w=3.8e-06 l=2e-06 c=5.2038e-14 as=2.31158e-13 ad=7.488e-13 ps=1.44e-06 pd=1.11673e-06 sim_w=2.88e-06 m_per_maxw=1.31944 numb_sub_cont=3 nfing=1 $X=-484300 $Y=276580 $D=21
M246 2 3 2 cpoly_p w=3.8e-06 l=2e-06 c=5.2038e-14 as=2.31158e-13 ad=7.488e-13 ps=1.44e-06 pd=1.11673e-06 sim_w=2.88e-06 m_per_maxw=1.31944 numb_sub_cont=3 nfing=1 $X=-481780 $Y=276580 $D=21
M247 2 3 2 cpoly_p w=3.8e-06 l=2e-06 c=5.2038e-14 as=2.31158e-13 ad=7.488e-13 ps=1.44e-06 pd=1.11673e-06 sim_w=2.88e-06 m_per_maxw=1.31944 numb_sub_cont=3 nfing=1 $X=-479260 $Y=276580 $D=21
M248 2 3 2 cpoly_p w=3.8e-06 l=2e-06 c=5.2038e-14 as=2.31158e-13 ad=7.488e-13 ps=1.44e-06 pd=1.11673e-06 sim_w=2.88e-06 m_per_maxw=1.31944 numb_sub_cont=3 nfing=1 $X=-476740 $Y=276580 $D=21
M249 2 3 2 cpoly_p w=3.8e-06 l=2e-06 c=5.2038e-14 as=2.31158e-13 ad=7.488e-13 ps=1.44e-06 pd=1.11673e-06 sim_w=2.88e-06 m_per_maxw=1.31944 numb_sub_cont=3 nfing=1 $X=-474220 $Y=276580 $D=21
M250 2 3 2 cpoly_p w=3.8e-06 l=2e-06 c=5.2038e-14 as=2.31158e-13 ad=7.488e-13 ps=1.44e-06 pd=1.11673e-06 sim_w=2.88e-06 m_per_maxw=1.31944 numb_sub_cont=3 nfing=1 $X=-471700 $Y=276580 $D=21
M251 2 3 2 cpoly_p w=3.8e-06 l=2e-06 c=5.2038e-14 as=2.31158e-13 ad=7.488e-13 ps=1.44e-06 pd=1.11673e-06 sim_w=2.88e-06 m_per_maxw=1.31944 numb_sub_cont=3 nfing=1 $X=-469180 $Y=276580 $D=21
M252 2 3 2 cpoly_p w=3.8e-06 l=2e-06 c=5.2038e-14 as=2.31158e-13 ad=7.488e-13 ps=1.44e-06 pd=1.11673e-06 sim_w=2.88e-06 m_per_maxw=1.31944 numb_sub_cont=3 nfing=1 $X=-466660 $Y=276580 $D=21
M253 2 3 2 cpoly_p w=3.8e-06 l=2e-06 c=5.2038e-14 as=2.31158e-13 ad=7.488e-13 ps=1.44e-06 pd=1.11673e-06 sim_w=2.88e-06 m_per_maxw=1.31944 numb_sub_cont=3 nfing=1 $X=-464140 $Y=276580 $D=21
M254 2 3 2 cpoly_p w=3.8e-06 l=2e-06 c=5.2038e-14 as=2.31158e-13 ad=7.488e-13 ps=1.44e-06 pd=1.11673e-06 sim_w=2.88e-06 m_per_maxw=1.31944 numb_sub_cont=3 nfing=1 $X=-461620 $Y=276580 $D=21
M255 2 3 2 cpoly_p w=3.8e-06 l=2e-06 c=5.2038e-14 as=2.31158e-13 ad=7.488e-13 ps=1.44e-06 pd=1.11673e-06 sim_w=2.88e-06 m_per_maxw=1.31944 numb_sub_cont=3 nfing=1 $X=-459100 $Y=276580 $D=21
M256 2 3 2 cpoly_p w=3.8e-06 l=2e-06 c=5.2038e-14 as=2.31158e-13 ad=7.488e-13 ps=1.44e-06 pd=1.11673e-06 sim_w=2.88e-06 m_per_maxw=1.31944 numb_sub_cont=3 nfing=1 $X=-456580 $Y=276580 $D=21
M257 2 3 2 cpoly_p w=3.8e-06 l=2e-06 c=5.2038e-14 as=2.31158e-13 ad=7.488e-13 ps=1.44e-06 pd=1.11673e-06 sim_w=2.88e-06 m_per_maxw=1.31944 numb_sub_cont=3 nfing=1 $X=-454060 $Y=276580 $D=21
M258 2 3 2 cpoly_p w=3.8e-06 l=2e-06 c=5.2038e-14 as=2.31158e-13 ad=7.488e-13 ps=1.44e-06 pd=1.11673e-06 sim_w=2.88e-06 m_per_maxw=1.31944 numb_sub_cont=3 nfing=1 $X=-451540 $Y=276580 $D=21
M259 2 3 2 cpoly_p w=3.8e-06 l=2e-06 c=5.2038e-14 as=2.31158e-13 ad=7.488e-13 ps=1.44e-06 pd=1.11673e-06 sim_w=2.88e-06 m_per_maxw=1.31944 numb_sub_cont=3 nfing=1 $X=-449020 $Y=276580 $D=21
M260 2 3 2 cpoly_p w=3.8e-06 l=2e-06 c=5.2038e-14 as=2.31158e-13 ad=7.488e-13 ps=1.44e-06 pd=1.11673e-06 sim_w=2.88e-06 m_per_maxw=1.31944 numb_sub_cont=3 nfing=1 $X=-446500 $Y=276580 $D=21
M261 2 3 2 cpoly_p w=3.8e-06 l=2e-06 c=5.2038e-14 as=2.31158e-13 ad=7.488e-13 ps=1.44e-06 pd=1.11673e-06 sim_w=2.88e-06 m_per_maxw=1.31944 numb_sub_cont=3 nfing=1 $X=-443980 $Y=276580 $D=21
M262 2 3 2 cpoly_p w=3.8e-06 l=2e-06 c=5.2038e-14 as=2.31158e-13 ad=7.488e-13 ps=1.44e-06 pd=1.11673e-06 sim_w=2.88e-06 m_per_maxw=1.31944 numb_sub_cont=3 nfing=1 $X=-441460 $Y=276580 $D=21
M263 2 3 2 cpoly_p w=3.8e-06 l=2e-06 c=5.2038e-14 as=2.31158e-13 ad=7.488e-13 ps=1.44e-06 pd=1.11673e-06 sim_w=2.88e-06 m_per_maxw=1.31944 numb_sub_cont=3 nfing=1 $X=-438940 $Y=276580 $D=21
M264 2 3 2 cpoly_p w=3.8e-06 l=2e-06 c=5.2038e-14 as=2.31158e-13 ad=7.488e-13 ps=1.44e-06 pd=1.11673e-06 sim_w=2.88e-06 m_per_maxw=1.31944 numb_sub_cont=3 nfing=1 $X=-436420 $Y=276580 $D=21
M265 2 3 2 cpoly_p w=3.8e-06 l=2e-06 c=5.2038e-14 as=2.31158e-13 ad=7.488e-13 ps=1.44e-06 pd=1.11673e-06 sim_w=2.88e-06 m_per_maxw=1.31944 numb_sub_cont=3 nfing=1 $X=-433900 $Y=276580 $D=21
M266 2 3 2 cpoly_p w=3.8e-06 l=2e-06 c=5.2038e-14 as=2.31158e-13 ad=7.488e-13 ps=1.44e-06 pd=1.11673e-06 sim_w=2.88e-06 m_per_maxw=1.31944 numb_sub_cont=3 nfing=1 $X=-431380 $Y=276580 $D=21
M267 2 3 2 cpoly_p w=3.8e-06 l=2e-06 c=5.2038e-14 as=2.31158e-13 ad=7.488e-13 ps=1.44e-06 pd=1.11673e-06 sim_w=2.88e-06 m_per_maxw=1.31944 numb_sub_cont=3 nfing=1 $X=-428860 $Y=276580 $D=21
M268 2 3 2 cpoly_p w=3.8e-06 l=2e-06 c=5.2038e-14 as=2.31158e-13 ad=7.488e-13 ps=1.44e-06 pd=1.11673e-06 sim_w=2.88e-06 m_per_maxw=1.31944 numb_sub_cont=3 nfing=1 $X=-426340 $Y=276580 $D=21
M269 2 3 2 cpoly_p w=3.8e-06 l=2e-06 c=5.2038e-14 as=2.31158e-13 ad=7.488e-13 ps=1.44e-06 pd=1.11673e-06 sim_w=2.88e-06 m_per_maxw=1.31944 numb_sub_cont=3 nfing=1 $X=-423820 $Y=276580 $D=21
M270 2 3 2 cpoly_p w=3.8e-06 l=2e-06 c=5.2038e-14 as=2.31158e-13 ad=7.488e-13 ps=1.44e-06 pd=1.11673e-06 sim_w=2.88e-06 m_per_maxw=1.31944 numb_sub_cont=3 nfing=1 $X=-421300 $Y=276580 $D=21
M271 2 3 2 cpoly_p w=3.8e-06 l=2e-06 c=5.2038e-14 as=2.31158e-13 ad=7.488e-13 ps=1.44e-06 pd=1.11673e-06 sim_w=2.88e-06 m_per_maxw=1.31944 numb_sub_cont=3 nfing=1 $X=-418780 $Y=276580 $D=21
M272 2 3 2 cpoly_p w=3.8e-06 l=2e-06 c=5.2038e-14 as=2.31158e-13 ad=7.488e-13 ps=1.44e-06 pd=1.11673e-06 sim_w=2.88e-06 m_per_maxw=1.31944 numb_sub_cont=3 nfing=1 $X=-416260 $Y=276580 $D=21
M273 2 3 2 cpoly_p w=3.8e-06 l=2e-06 c=5.2038e-14 as=2.31158e-13 ad=7.488e-13 ps=1.44e-06 pd=1.11673e-06 sim_w=2.88e-06 m_per_maxw=1.31944 numb_sub_cont=3 nfing=1 $X=-413740 $Y=276580 $D=21
M274 2 3 2 cpoly_p w=3.8e-06 l=2e-06 c=5.2038e-14 as=2.31158e-13 ad=7.488e-13 ps=1.44e-06 pd=1.11673e-06 sim_w=2.88e-06 m_per_maxw=1.31944 numb_sub_cont=3 nfing=1 $X=-411220 $Y=276580 $D=21
M275 2 3 2 cpoly_p w=3.8e-06 l=2e-06 c=5.2038e-14 as=2.31158e-13 ad=7.488e-13 ps=1.44e-06 pd=1.11673e-06 sim_w=2.88e-06 m_per_maxw=1.31944 numb_sub_cont=3 nfing=1 $X=-408700 $Y=276580 $D=21
M276 2 3 2 cpoly_p w=3.8e-06 l=2e-06 c=5.2038e-14 as=2.31158e-13 ad=7.488e-13 ps=1.44e-06 pd=1.11673e-06 sim_w=2.88e-06 m_per_maxw=1.31944 numb_sub_cont=3 nfing=1 $X=-406180 $Y=276580 $D=21
M277 2 3 2 cpoly_p w=3.8e-06 l=2e-06 c=5.2038e-14 as=2.31158e-13 ad=7.488e-13 ps=1.44e-06 pd=1.11673e-06 sim_w=2.88e-06 m_per_maxw=1.31944 numb_sub_cont=3 nfing=1 $X=-403660 $Y=276580 $D=21
M278 2 3 2 cpoly_p w=3.8e-06 l=2e-06 c=5.2038e-14 as=2.31158e-13 ad=7.488e-13 ps=1.44e-06 pd=1.11673e-06 sim_w=2.88e-06 m_per_maxw=1.31944 numb_sub_cont=3 nfing=1 $X=-401140 $Y=276580 $D=21
M279 3 2 3 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=1.67141e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=-1013280 $Y=283540 $D=22
M280 3 2 3 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=-1010760 $Y=283540 $D=22
M281 3 2 3 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=-1008240 $Y=283540 $D=22
M282 3 2 3 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=-1005720 $Y=283540 $D=22
M283 3 2 3 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=-1003200 $Y=283540 $D=22
M284 3 2 3 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=-1000680 $Y=283540 $D=22
M285 3 2 3 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=-998160 $Y=283540 $D=22
M286 3 2 3 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=-995640 $Y=283540 $D=22
M287 3 2 3 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=-993120 $Y=283540 $D=22
M288 3 2 3 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=-990600 $Y=283540 $D=22
M289 3 2 3 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=-988080 $Y=283540 $D=22
M290 3 2 3 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=-985560 $Y=283540 $D=22
M291 3 2 3 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=-983040 $Y=283540 $D=22
M292 3 2 3 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=-980520 $Y=283540 $D=22
M293 3 2 3 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=-978000 $Y=283540 $D=22
M294 3 2 3 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=-975480 $Y=283540 $D=22
M295 3 2 3 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=-972960 $Y=283540 $D=22
M296 3 2 3 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=-970440 $Y=283540 $D=22
M297 3 2 3 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=-967920 $Y=283540 $D=22
M298 3 2 3 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=-965400 $Y=283540 $D=22
M299 3 2 3 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=-962880 $Y=283540 $D=22
M300 3 2 3 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=-960360 $Y=283540 $D=22
M301 3 2 3 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=-957840 $Y=283540 $D=22
M302 3 2 3 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=-955320 $Y=283540 $D=22
M303 3 2 3 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=-952800 $Y=283540 $D=22
M304 3 2 3 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=-950280 $Y=283540 $D=22
M305 3 2 3 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=-947760 $Y=283540 $D=22
M306 3 2 3 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=-945240 $Y=283540 $D=22
M307 3 2 3 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=-942720 $Y=283540 $D=22
M308 3 2 3 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=-940200 $Y=283540 $D=22
M309 3 2 3 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=-937680 $Y=283540 $D=22
M310 3 2 3 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=-935160 $Y=283540 $D=22
M311 3 2 3 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=-932640 $Y=283540 $D=22
M312 3 2 3 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=-930120 $Y=283540 $D=22
M313 3 2 3 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=-927600 $Y=283540 $D=22
M314 3 2 3 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=-925080 $Y=283540 $D=22
M315 3 2 3 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=-922560 $Y=283540 $D=22
M316 3 2 3 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=-920040 $Y=283540 $D=22
M317 3 2 3 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=-917520 $Y=283540 $D=22
M318 3 2 3 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=-915000 $Y=283540 $D=22
M319 3 2 3 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=-912480 $Y=283540 $D=22
M320 3 2 3 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=-909960 $Y=283540 $D=22
M321 3 2 3 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=-907440 $Y=283540 $D=22
M322 3 2 3 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=-904920 $Y=283540 $D=22
M323 3 2 3 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=-902400 $Y=283540 $D=22
M324 3 2 3 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=-899880 $Y=283540 $D=22
M325 3 2 3 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=-897360 $Y=283540 $D=22
M326 3 2 3 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=-894840 $Y=283540 $D=22
M327 3 2 3 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=-892320 $Y=283540 $D=22
M328 3 2 3 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=-889800 $Y=283540 $D=22
M329 3 2 3 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=-887280 $Y=283540 $D=22
M330 3 2 3 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=-884760 $Y=283540 $D=22
M331 3 2 3 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=-882240 $Y=283540 $D=22
M332 3 2 3 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=-879720 $Y=283540 $D=22
M333 3 2 3 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=-877200 $Y=283540 $D=22
M334 3 2 3 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=-874680 $Y=283540 $D=22
M335 3 2 3 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=-872160 $Y=283540 $D=22
M336 3 2 3 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=-869640 $Y=283540 $D=22
M337 3 2 3 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=-867120 $Y=283540 $D=22
M338 3 2 3 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=-864600 $Y=283540 $D=22
M339 3 2 3 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=-862080 $Y=283540 $D=22
M340 3 2 3 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=-859560 $Y=283540 $D=22
M341 3 2 3 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=-857040 $Y=283540 $D=22
M342 3 2 3 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=-854520 $Y=283540 $D=22
M343 3 2 3 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=-852000 $Y=283540 $D=22
M344 3 2 3 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=-849480 $Y=283540 $D=22
M345 3 2 3 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=-846960 $Y=283540 $D=22
M346 3 2 3 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=-844440 $Y=283540 $D=22
M347 3 2 3 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=-841920 $Y=283540 $D=22
M348 3 2 3 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=-839400 $Y=283540 $D=22
M349 3 2 3 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=-836880 $Y=283540 $D=22
M350 3 2 3 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=-834360 $Y=283540 $D=22
M351 3 2 3 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=-831840 $Y=283540 $D=22
M352 3 2 3 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=-829320 $Y=283540 $D=22
M353 3 2 3 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=-826800 $Y=283540 $D=22
M354 3 2 3 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=-824280 $Y=283540 $D=22
M355 3 2 3 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=-821760 $Y=283540 $D=22
M356 3 2 3 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=-819240 $Y=283540 $D=22
M357 3 2 3 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=-816720 $Y=283540 $D=22
M358 3 2 3 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=-814200 $Y=283540 $D=22
M359 3 2 3 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=-811680 $Y=283540 $D=22
M360 3 2 3 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=-809160 $Y=283540 $D=22
M361 3 2 3 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=-806640 $Y=283540 $D=22
M362 3 2 3 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=-804120 $Y=283540 $D=22
M363 3 2 3 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=-801600 $Y=283540 $D=22
M364 3 2 3 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=-799080 $Y=283540 $D=22
M365 3 2 3 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=-796560 $Y=283540 $D=22
M366 3 2 3 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=-794040 $Y=283540 $D=22
M367 3 2 3 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=-791520 $Y=283540 $D=22
M368 3 2 3 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=-789000 $Y=283540 $D=22
M369 3 2 3 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=-786480 $Y=283540 $D=22
M370 3 2 3 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=-783960 $Y=283540 $D=22
M371 3 2 3 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=-781440 $Y=283540 $D=22
M372 3 2 3 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=-778920 $Y=283540 $D=22
M373 3 2 3 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=-776400 $Y=283540 $D=22
M374 3 2 3 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=-773880 $Y=283540 $D=22
M375 3 2 3 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=-771360 $Y=283540 $D=22
M376 3 2 3 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=-768840 $Y=283540 $D=22
M377 3 2 3 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=-766320 $Y=283540 $D=22
M378 3 2 3 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=-763800 $Y=283540 $D=22
M379 3 2 3 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=-761280 $Y=283540 $D=22
M380 3 2 3 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=-758760 $Y=283540 $D=22
M381 3 2 3 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=-756240 $Y=283540 $D=22
M382 3 2 3 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=-753720 $Y=283540 $D=22
M383 3 2 3 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=-751200 $Y=283540 $D=22
M384 3 2 3 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=-748680 $Y=283540 $D=22
M385 3 2 3 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=-746160 $Y=283540 $D=22
M386 3 2 3 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=-743640 $Y=283540 $D=22
M387 3 2 3 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=-741120 $Y=283540 $D=22
M388 3 2 3 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=-738600 $Y=283540 $D=22
M389 3 2 3 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=-736080 $Y=283540 $D=22
M390 3 2 3 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=-733560 $Y=283540 $D=22
M391 3 2 3 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=-731040 $Y=283540 $D=22
M392 3 2 3 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=-728520 $Y=283540 $D=22
M393 3 2 3 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=-726000 $Y=283540 $D=22
M394 3 2 3 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=-723480 $Y=283540 $D=22
M395 3 2 3 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=-720960 $Y=283540 $D=22
M396 3 2 3 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=-718440 $Y=283540 $D=22
M397 3 2 3 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=-715920 $Y=283540 $D=22
M398 3 2 3 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=-713400 $Y=283540 $D=22
M399 3 2 3 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=-710880 $Y=283540 $D=22
M400 3 2 3 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=-708360 $Y=283540 $D=22
M401 3 2 3 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=-705840 $Y=283540 $D=22
M402 3 2 3 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=-703320 $Y=283540 $D=22
M403 3 2 3 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=-700800 $Y=283540 $D=22
M404 3 2 3 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=-698280 $Y=283540 $D=22
M405 3 2 3 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=-695760 $Y=283540 $D=22
M406 3 2 3 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=-693240 $Y=283540 $D=22
M407 3 2 3 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=-690720 $Y=283540 $D=22
M408 3 2 3 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=-688200 $Y=283540 $D=22
M409 3 2 3 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=-685680 $Y=283540 $D=22
M410 3 2 3 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=-683160 $Y=283540 $D=22
M411 3 2 3 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=-680640 $Y=283540 $D=22
M412 3 2 3 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=-678120 $Y=283540 $D=22
M413 3 2 3 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=-675600 $Y=283540 $D=22
M414 3 2 3 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=-673080 $Y=283540 $D=22
M415 3 2 3 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=-670560 $Y=283540 $D=22
M416 3 2 3 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=-668040 $Y=283540 $D=22
M417 3 2 3 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=-665520 $Y=283540 $D=22
M418 3 2 3 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=-663000 $Y=283540 $D=22
M419 3 2 3 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=-660480 $Y=283540 $D=22
M420 3 2 3 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=-657960 $Y=283540 $D=22
M421 3 2 3 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=-655440 $Y=283540 $D=22
M422 3 2 3 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=-652920 $Y=283540 $D=22
M423 3 2 3 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=-650400 $Y=283540 $D=22
M424 3 2 3 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=-647880 $Y=283540 $D=22
M425 3 2 3 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=-645360 $Y=283540 $D=22
M426 3 2 3 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=-642840 $Y=283540 $D=22
M427 3 2 3 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=-640320 $Y=283540 $D=22
M428 3 2 3 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=-637800 $Y=283540 $D=22
M429 3 2 3 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=-635280 $Y=283540 $D=22
M430 3 2 3 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=-632760 $Y=283540 $D=22
M431 3 2 3 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=-630240 $Y=283540 $D=22
M432 3 2 3 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=-627720 $Y=283540 $D=22
M433 3 2 3 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=-625200 $Y=283540 $D=22
M434 3 2 3 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=-622680 $Y=283540 $D=22
M435 3 2 3 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=-620160 $Y=283540 $D=22
M436 3 2 3 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=-617640 $Y=283540 $D=22
M437 3 2 3 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=-615120 $Y=283540 $D=22
M438 3 2 3 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=-612600 $Y=283540 $D=22
M439 3 2 3 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=-610080 $Y=283540 $D=22
M440 3 2 3 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=-607560 $Y=283540 $D=22
M441 3 2 3 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=-605040 $Y=283540 $D=22
M442 3 2 3 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=-602520 $Y=283540 $D=22
M443 3 2 3 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=-600000 $Y=283540 $D=22
M444 3 2 3 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=-597480 $Y=283540 $D=22
M445 3 2 3 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=-594960 $Y=283540 $D=22
M446 3 2 3 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=-592440 $Y=283540 $D=22
M447 3 2 3 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=-589920 $Y=283540 $D=22
M448 3 2 3 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=-587400 $Y=283540 $D=22
M449 3 2 3 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=-584880 $Y=283540 $D=22
M450 3 2 3 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=-582360 $Y=283540 $D=22
M451 3 2 3 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=-579840 $Y=283540 $D=22
M452 3 2 3 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=-577320 $Y=283540 $D=22
M453 3 2 3 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=-574800 $Y=283540 $D=22
M454 3 2 3 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=-572280 $Y=283540 $D=22
M455 3 2 3 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=-569760 $Y=283540 $D=22
M456 3 2 3 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=-567240 $Y=283540 $D=22
M457 3 2 3 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=-564720 $Y=283540 $D=22
M458 3 2 3 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=-562200 $Y=283540 $D=22
M459 3 2 3 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=-559680 $Y=283540 $D=22
M460 3 2 3 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=-557160 $Y=283540 $D=22
M461 3 2 3 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=-554640 $Y=283540 $D=22
M462 3 2 3 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=-552120 $Y=283540 $D=22
M463 3 2 3 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=-549600 $Y=283540 $D=22
M464 3 2 3 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=-547080 $Y=283540 $D=22
M465 3 2 3 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=-544560 $Y=283540 $D=22
M466 3 2 3 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=-542040 $Y=283540 $D=22
M467 3 2 3 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=-539520 $Y=283540 $D=22
M468 3 2 3 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=-537000 $Y=283540 $D=22
M469 3 2 3 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=-534480 $Y=283540 $D=22
M470 3 2 3 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=-531960 $Y=283540 $D=22
M471 3 2 3 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=-529440 $Y=283540 $D=22
M472 3 2 3 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=-526920 $Y=283540 $D=22
M473 3 2 3 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=-524400 $Y=283540 $D=22
M474 3 2 3 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=-521880 $Y=283540 $D=22
M475 3 2 3 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=-519360 $Y=283540 $D=22
M476 3 2 3 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=-516840 $Y=283540 $D=22
M477 3 2 3 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=-514320 $Y=283540 $D=22
M478 3 2 3 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=-511800 $Y=283540 $D=22
M479 3 2 3 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=-509280 $Y=283540 $D=22
M480 3 2 3 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=-506760 $Y=283540 $D=22
M481 3 2 3 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=-504240 $Y=283540 $D=22
M482 3 2 3 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=-501720 $Y=283540 $D=22
M483 3 2 3 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=-499200 $Y=283540 $D=22
M484 3 2 3 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=-496680 $Y=283540 $D=22
M485 3 2 3 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=-494160 $Y=283540 $D=22
M486 3 2 3 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=-491640 $Y=283540 $D=22
M487 3 2 3 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=-489120 $Y=283540 $D=22
M488 3 2 3 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=-486600 $Y=283540 $D=22
M489 3 2 3 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=-484080 $Y=283540 $D=22
M490 3 2 3 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=-481560 $Y=283540 $D=22
M491 3 2 3 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=-479040 $Y=283540 $D=22
M492 3 2 3 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=-476520 $Y=283540 $D=22
M493 3 2 3 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=-474000 $Y=283540 $D=22
M494 3 2 3 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=-471480 $Y=283540 $D=22
M495 3 2 3 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=-468960 $Y=283540 $D=22
M496 3 2 3 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=-466440 $Y=283540 $D=22
M497 3 2 3 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=-463920 $Y=283540 $D=22
M498 3 2 3 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=-461400 $Y=283540 $D=22
M499 3 2 3 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=-458880 $Y=283540 $D=22
M500 3 2 3 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=-456360 $Y=283540 $D=22
M501 3 2 3 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=-453840 $Y=283540 $D=22
M502 3 2 3 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=-451320 $Y=283540 $D=22
M503 3 2 3 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=-448800 $Y=283540 $D=22
M504 3 2 3 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=-446280 $Y=283540 $D=22
M505 3 2 3 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=-443760 $Y=283540 $D=22
M506 3 2 3 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=-441240 $Y=283540 $D=22
M507 3 2 3 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=-438720 $Y=283540 $D=22
M508 3 2 3 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=-436200 $Y=283540 $D=22
M509 3 2 3 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=-433680 $Y=283540 $D=22
M510 3 2 3 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=-431160 $Y=283540 $D=22
M511 3 2 3 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=-428640 $Y=283540 $D=22
M512 3 2 3 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=-426120 $Y=283540 $D=22
M513 3 2 3 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=-423600 $Y=283540 $D=22
M514 3 2 3 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=-421080 $Y=283540 $D=22
M515 3 2 3 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=-418560 $Y=283540 $D=22
M516 3 2 3 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=-416040 $Y=283540 $D=22
M517 3 2 3 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=-413520 $Y=283540 $D=22
M518 3 2 3 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=-411000 $Y=283540 $D=22
M519 3 2 3 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=-408480 $Y=283540 $D=22
M520 3 2 3 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=-405960 $Y=283540 $D=22
M521 3 2 3 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=-403440 $Y=283540 $D=22
M522 3 2 3 cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=-400920 $Y=283540 $D=22
X523 3 16 13 pmos_a_CDNS_5887047866540 $T=-1007680 272760 1 0 $X=-1007680 $Y=270560
X525 14 15 17 16 Cell_Usub $T=-401880 271760 1 0 $X=-402240 $Y=268540
X526 14 15 17 16 Cell_Usub $T=-401880 271760 0 0 $X=-402240 $Y=271420
X527 14 15 17 16 ICV_158 $T=-426040 271760 1 0 $X=-426400 $Y=268540
X528 14 15 17 16 ICV_159 $T=-1005880 271760 1 0 $X=-1006240 $Y=268540
X529 14 15 17 16 ICV_159 $T=-957560 271760 1 0 $X=-957920 $Y=268540
X530 14 15 17 16 ICV_159 $T=-909240 271760 1 0 $X=-909600 $Y=268540
X531 14 15 17 16 ICV_159 $T=-860920 271760 1 0 $X=-861280 $Y=268540
X532 14 15 17 16 ICV_159 $T=-812600 271760 1 0 $X=-812960 $Y=268540
X533 14 15 17 16 ICV_159 $T=-764280 271760 1 0 $X=-764640 $Y=268540
X534 14 15 17 16 ICV_159 $T=-715960 271760 1 0 $X=-716320 $Y=268540
X535 14 15 17 16 ICV_159 $T=-667640 271760 1 0 $X=-668000 $Y=268540
X536 14 15 17 16 ICV_159 $T=-619320 271760 1 0 $X=-619680 $Y=268540
X537 14 15 17 16 ICV_159 $T=-571000 271760 1 0 $X=-571360 $Y=268540
X538 14 15 17 16 ICV_159 $T=-522680 271760 1 0 $X=-523040 $Y=268540
X539 14 15 17 16 ICV_159 $T=-474360 271760 1 0 $X=-474720 $Y=268540
.ENDS
***************************************
.SUBCKT ICV_161
** N=5 EP=0 IP=0 FDC=0
*.SEEDPROM
.ENDS
***************************************
.SUBCKT ICV_162
** N=2 EP=0 IP=0 FDC=0
*.SEEDPROM
.ENDS
***************************************
.SUBCKT nmos_a_CDNS_5887047866548
** N=3 EP=0 IP=0 FDC=0
*.SEEDPROM
.ENDS
***************************************
.SUBCKT ICV_163 5 6 7
** N=9 EP=3 IP=3 FDC=1
*.SEEDPROM
M0 7 6 5 5 nmos_a L=2.8e-07 W=4.2e-06 AD=1.59086e-12 AS=1.68e-12 PD=3.97714e-06 PS=1.98857e-06 w_cont=1.6e-06 nfing=1 source_num=2 $X=-436680 $Y=-35320 $D=1
.ENDS
***************************************
.SUBCKT dn_CDNS_5887047866549 1 2
** N=2 EP=2 IP=0 FDC=1
D0 2 1 dn PJ=2e-05 m=1 $X=-460 $Y=0 $D=9
.ENDS
***************************************
.SUBCKT ICV_164 3 4 7 8
** N=11 EP=4 IP=13 FDC=6
*.SEEDPROM
M0 8 4 3 3 nmos_a L=2.8e-07 W=4.2e-06 AD=1.59086e-12 AS=2.23341e-12 PD=3.97714e-06 PS=1.98857e-06 w_cont=1.6e-06 nfing=1 source_num=2 $X=-436840 $Y=-42920 $D=1
X2 3 7 dn_CDNS_5887047866549 $T=-436660 -146660 0 0 $X=-437300 $Y=-146960
X3 7 9 dn_CDNS_5887047866549 $T=-436660 -126060 0 0 $X=-437300 $Y=-126360
X4 9 10 dn_CDNS_5887047866549 $T=-436660 -105460 0 0 $X=-437300 $Y=-105760
X5 10 11 dn_CDNS_5887047866549 $T=-436660 -84860 0 0 $X=-437300 $Y=-85160
X6 11 4 dn_CDNS_5887047866549 $T=-436660 -64260 0 0 $X=-437300 $Y=-64560
.ENDS
***************************************
.SUBCKT ICV_165
** N=41 EP=0 IP=0 FDC=0
*.SEEDPROM
.ENDS
***************************************
.SUBCKT dn_CDNS_5887047866561
** N=2 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT Usub_7V gnd! vdd! nTest Usub
** N=58 EP=4 IP=621 FDC=4091
M0 gnd! 21 gnd! gnd! nmos_a L=2e-06 W=5.5e-06 AD=8.30487e-13 AS=1.43e-12 PD=1.59709e-06 PS=1.59709e-06 w_cont=6e-07 nfing=1 source_num=2 $X=-196340 $Y=275380 $D=1
M1 vdd! gnd! vdd! vdd! nmos_a L=2e-06 W=6.5e-06 AD=8.1792e-13 AS=2.6e-12 PD=1.57292e-06 PS=1.57292e-06 w_cont=6e-07 nfing=1 source_num=2 $X=-182520 $Y=265080 $D=1
M2 vdd! gnd! vdd! vdd! nmos_a L=2e-06 W=6.5e-06 AD=8.1792e-13 AS=3.38e-12 PD=1.57292e-06 PS=1.57292e-06 w_cont=6e-07 nfing=1 source_num=2 $X=-180000 $Y=265080 $D=1
M3 vdd! gnd! vdd! vdd! nmos_a L=2e-06 W=6.5e-06 AD=8.1792e-13 AS=3.38e-12 PD=1.57292e-06 PS=1.57292e-06 w_cont=6e-07 nfing=1 source_num=2 $X=-177480 $Y=265080 $D=1
M4 vdd! gnd! vdd! vdd! nmos_a L=2e-06 W=6.5e-06 AD=8.1792e-13 AS=3.38e-12 PD=1.57292e-06 PS=1.57292e-06 w_cont=6e-07 nfing=1 source_num=2 $X=-174960 $Y=265080 $D=1
M5 vdd! gnd! vdd! vdd! nmos_a L=2e-06 W=6.5e-06 AD=8.1792e-13 AS=3.38e-12 PD=1.57292e-06 PS=1.57292e-06 w_cont=6e-07 nfing=1 source_num=2 $X=-172440 $Y=265080 $D=1
M6 vdd! gnd! vdd! vdd! nmos_a L=2e-06 W=6.5e-06 AD=8.1792e-13 AS=3.38e-12 PD=1.57292e-06 PS=1.57292e-06 w_cont=6e-07 nfing=1 source_num=2 $X=-169920 $Y=265080 $D=1
M7 vdd! gnd! vdd! vdd! nmos_a L=2e-06 W=6.5e-06 AD=8.1792e-13 AS=3.38e-12 PD=1.57292e-06 PS=1.57292e-06 w_cont=6e-07 nfing=1 source_num=2 $X=-167400 $Y=265080 $D=1
M8 vdd! gnd! vdd! vdd! nmos_a L=2e-06 W=6.5e-06 AD=8.1792e-13 AS=3.38e-12 PD=1.57292e-06 PS=1.57292e-06 w_cont=6e-07 nfing=1 source_num=2 $X=-164880 $Y=265080 $D=1
M9 vdd! gnd! vdd! vdd! nmos_a L=2e-06 W=6.5e-06 AD=8.1792e-13 AS=3.38e-12 PD=1.57292e-06 PS=1.57292e-06 w_cont=6e-07 nfing=1 source_num=2 $X=-162360 $Y=265080 $D=1
M10 vdd! gnd! vdd! vdd! nmos_a L=2e-06 W=6.5e-06 AD=8.1792e-13 AS=3.38e-12 PD=1.57292e-06 PS=1.57292e-06 w_cont=6e-07 nfing=1 source_num=2 $X=-159840 $Y=265080 $D=1
M11 vdd! gnd! vdd! vdd! nmos_a L=2e-06 W=6.5e-06 AD=8.1792e-13 AS=3.38e-12 PD=1.57292e-06 PS=1.57292e-06 w_cont=6e-07 nfing=1 source_num=2 $X=-157320 $Y=265080 $D=1
M12 vdd! gnd! vdd! vdd! nmos_a L=2e-06 W=6.5e-06 AD=8.1792e-13 AS=3.38e-12 PD=1.57292e-06 PS=1.57292e-06 w_cont=6e-07 nfing=1 source_num=2 $X=-154800 $Y=265080 $D=1
M13 vdd! gnd! vdd! vdd! nmos_a L=2e-06 W=6.5e-06 AD=8.1792e-13 AS=3.38e-12 PD=1.57292e-06 PS=1.57292e-06 w_cont=6e-07 nfing=1 source_num=2 $X=-152280 $Y=265080 $D=1
M14 vdd! gnd! vdd! vdd! nmos_a L=2e-06 W=6.5e-06 AD=8.1792e-13 AS=3.38e-12 PD=1.57292e-06 PS=1.57292e-06 w_cont=6e-07 nfing=1 source_num=2 $X=-149760 $Y=265080 $D=1
M15 vdd! gnd! vdd! vdd! nmos_a L=2e-06 W=6.5e-06 AD=8.1792e-13 AS=3.38e-12 PD=1.57292e-06 PS=1.57292e-06 w_cont=6e-07 nfing=1 source_num=2 $X=-147240 $Y=265080 $D=1
M16 vdd! gnd! vdd! vdd! nmos_a L=2e-06 W=6.5e-06 AD=8.1792e-13 AS=3.38e-12 PD=1.57292e-06 PS=1.57292e-06 w_cont=6e-07 nfing=1 source_num=2 $X=-144720 $Y=265080 $D=1
M17 vdd! gnd! vdd! vdd! nmos_a L=2e-06 W=6.5e-06 AD=8.1792e-13 AS=3.38e-12 PD=1.57292e-06 PS=1.57292e-06 w_cont=6e-07 nfing=1 source_num=2 $X=-142200 $Y=265080 $D=1
M18 vdd! gnd! vdd! vdd! nmos_a L=2e-06 W=6.5e-06 AD=8.1792e-13 AS=3.38e-12 PD=1.57292e-06 PS=1.57292e-06 w_cont=6e-07 nfing=1 source_num=2 $X=-139680 $Y=265080 $D=1
M19 vdd! gnd! vdd! vdd! nmos_a L=2e-06 W=6.5e-06 AD=8.1792e-13 AS=3.38e-12 PD=1.57292e-06 PS=1.57292e-06 w_cont=6e-07 nfing=1 source_num=2 $X=-137160 $Y=265080 $D=1
M20 vdd! gnd! vdd! vdd! nmos_a L=2e-06 W=6.5e-06 AD=8.1792e-13 AS=3.38e-12 PD=1.57292e-06 PS=1.57292e-06 w_cont=6e-07 nfing=1 source_num=2 $X=-134640 $Y=265080 $D=1
M21 vdd! gnd! vdd! vdd! nmos_a L=2e-06 W=6.5e-06 AD=8.1792e-13 AS=3.38e-12 PD=1.57292e-06 PS=1.57292e-06 w_cont=6e-07 nfing=1 source_num=2 $X=-132120 $Y=265080 $D=1
M22 vdd! gnd! vdd! vdd! nmos_a L=2e-06 W=6.5e-06 AD=8.1792e-13 AS=3.38e-12 PD=1.57292e-06 PS=1.57292e-06 w_cont=6e-07 nfing=1 source_num=2 $X=-129600 $Y=265080 $D=1
M23 vdd! gnd! vdd! vdd! nmos_a L=2e-06 W=6.5e-06 AD=8.1792e-13 AS=3.38e-12 PD=1.57292e-06 PS=1.57292e-06 w_cont=6e-07 nfing=1 source_num=2 $X=-127080 $Y=265080 $D=1
M24 vdd! gnd! vdd! vdd! nmos_a L=2e-06 W=6.5e-06 AD=8.1792e-13 AS=3.38e-12 PD=1.57292e-06 PS=1.57292e-06 w_cont=6e-07 nfing=1 source_num=2 $X=-124560 $Y=265080 $D=1
M25 vdd! gnd! vdd! vdd! nmos_a L=2e-06 W=6.5e-06 AD=8.1792e-13 AS=3.38e-12 PD=1.57292e-06 PS=1.57292e-06 w_cont=6e-07 nfing=1 source_num=2 $X=-122040 $Y=265080 $D=1
M26 vdd! gnd! vdd! vdd! nmos_a L=2e-06 W=6.5e-06 AD=8.1792e-13 AS=3.38e-12 PD=1.57292e-06 PS=1.57292e-06 w_cont=6e-07 nfing=1 source_num=2 $X=-119520 $Y=265080 $D=1
M27 vdd! gnd! vdd! vdd! nmos_a L=2e-06 W=6.5e-06 AD=8.1792e-13 AS=3.38e-12 PD=1.57292e-06 PS=1.57292e-06 w_cont=6e-07 nfing=1 source_num=2 $X=-117000 $Y=265080 $D=1
M28 vdd! gnd! vdd! vdd! nmos_a L=2e-06 W=6.5e-06 AD=8.1792e-13 AS=3.38e-12 PD=1.57292e-06 PS=1.57292e-06 w_cont=6e-07 nfing=1 source_num=2 $X=-114480 $Y=265080 $D=1
M29 vdd! gnd! vdd! vdd! nmos_a L=2e-06 W=6.5e-06 AD=8.1792e-13 AS=3.38e-12 PD=1.57292e-06 PS=1.57292e-06 w_cont=6e-07 nfing=1 source_num=2 $X=-111960 $Y=265080 $D=1
M30 vdd! gnd! vdd! vdd! nmos_a L=2e-06 W=6.5e-06 AD=8.1792e-13 AS=3.38e-12 PD=1.57292e-06 PS=1.57292e-06 w_cont=6e-07 nfing=1 source_num=2 $X=-109440 $Y=265080 $D=1
M31 vdd! gnd! vdd! vdd! nmos_a L=2e-06 W=6.5e-06 AD=8.1792e-13 AS=3.38e-12 PD=1.57292e-06 PS=1.57292e-06 w_cont=6e-07 nfing=1 source_num=2 $X=-106920 $Y=265080 $D=1
M32 vdd! gnd! vdd! vdd! nmos_a L=2e-06 W=6.5e-06 AD=8.1792e-13 AS=3.38e-12 PD=1.57292e-06 PS=1.57292e-06 w_cont=6e-07 nfing=1 source_num=2 $X=-104400 $Y=265080 $D=1
M33 vdd! gnd! vdd! vdd! nmos_a L=2e-06 W=6.5e-06 AD=8.1792e-13 AS=3.38e-12 PD=1.57292e-06 PS=1.57292e-06 w_cont=6e-07 nfing=1 source_num=2 $X=-101880 $Y=265080 $D=1
M34 vdd! gnd! vdd! vdd! nmos_a L=2e-06 W=6.5e-06 AD=8.1792e-13 AS=3.38e-12 PD=1.57292e-06 PS=1.57292e-06 w_cont=6e-07 nfing=1 source_num=2 $X=-99360 $Y=265080 $D=1
M35 vdd! gnd! vdd! vdd! nmos_a L=2e-06 W=6.5e-06 AD=8.1792e-13 AS=3.38e-12 PD=1.57292e-06 PS=1.57292e-06 w_cont=6e-07 nfing=1 source_num=2 $X=-96840 $Y=265080 $D=1
M36 vdd! gnd! vdd! vdd! nmos_a L=2e-06 W=6.5e-06 AD=8.1792e-13 AS=3.38e-12 PD=1.57292e-06 PS=1.57292e-06 w_cont=6e-07 nfing=1 source_num=2 $X=-94320 $Y=265080 $D=1
M37 vdd! gnd! vdd! vdd! nmos_a L=2e-06 W=6.5e-06 AD=8.1792e-13 AS=3.38e-12 PD=1.57292e-06 PS=1.57292e-06 w_cont=6e-07 nfing=1 source_num=2 $X=-91800 $Y=265080 $D=1
M38 vdd! gnd! vdd! vdd! nmos_a L=2e-06 W=6.5e-06 AD=8.1792e-13 AS=3.38e-12 PD=1.57292e-06 PS=1.57292e-06 w_cont=6e-07 nfing=1 source_num=2 $X=-89280 $Y=265080 $D=1
M39 vdd! gnd! vdd! vdd! nmos_a L=2e-06 W=6.5e-06 AD=8.1792e-13 AS=3.38e-12 PD=1.57292e-06 PS=1.57292e-06 w_cont=6e-07 nfing=1 source_num=2 $X=-86760 $Y=265080 $D=1
M40 vdd! gnd! vdd! vdd! nmos_a L=2e-06 W=6.5e-06 AD=8.1792e-13 AS=2.6e-12 PD=1.57292e-06 PS=1.57292e-06 w_cont=6e-07 nfing=1 source_num=2 $X=-84240 $Y=265080 $D=1
M41 24 45 vdd! vdd! pmos_a L=2.4e-07 W=5e-07 AD=4.4e-13 AS=1.585e-13 PD=1.1e-06 PS=5.5e-07 w_cont=6e-07 nfing=1 mmm=1 $X=-195580 $Y=267740 $D=5
M42 24 26 vdd! vdd! pmos_a L=2.4e-07 W=5e-07 AD=4.4e-13 AS=1.585e-13 PD=1.1e-06 PS=5.5e-07 w_cont=6e-07 nfing=1 mmm=1 $X=-194820 $Y=267740 $D=5
M43 26 24 vdd! vdd! pmos_a L=2.4e-07 W=5e-07 AD=4.4e-13 AS=1.585e-13 PD=1.1e-06 PS=5.5e-07 w_cont=6e-07 nfing=1 mmm=1 $X=-193400 $Y=267740 $D=5
M44 26 27 vdd! vdd! pmos_a L=2.4e-07 W=5e-07 AD=4.4e-13 AS=1.585e-13 PD=1.1e-06 PS=5.5e-07 w_cont=6e-07 nfing=1 mmm=1 $X=-192640 $Y=267740 $D=5
M45 27 53 49 49 pmos_a L=2.4e-07 W=4.8e-07 AD=4.32e-13 AS=1.224e-13 PD=1.08e-06 PS=5.4e-07 w_cont=6e-07 nfing=1 mmm=1 $X=-190960 $Y=267620 $D=5
M46 29 26 vdd! vdd! pmos_a L=2.4e-07 W=2.6e-06 AD=1.28e-12 AS=1.69e-13 PD=3.2e-06 PS=1.6e-06 w_cont=6e-07 nfing=1 mmm=1 $X=-185300 $Y=267660 $D=5
M47 29 26 vdd! vdd! pmos_a L=2.4e-07 W=2.6e-06 AD=1.28e-12 AS=1.69e-13 PD=3.2e-06 PS=1.6e-06 w_cont=6e-07 nfing=1 mmm=1 $X=-184540 $Y=267660 $D=5
M48 43 24 vdd! vdd! pmos_a L=2.4e-07 W=2.6e-06 AD=1.28e-12 AS=1.69e-13 PD=3.2e-06 PS=1.6e-06 w_cont=6e-07 nfing=1 mmm=1 $X=-203700 $Y=267660 $D=5
M49 43 24 vdd! vdd! pmos_a L=2.4e-07 W=2.6e-06 AD=1.28e-12 AS=1.69e-13 PD=3.2e-06 PS=1.6e-06 w_cont=6e-07 nfing=1 mmm=1 $X=-202940 $Y=267660 $D=5
M50 45 56 51 51 pmos_a L=2.4e-07 W=4.8e-07 AD=4.32e-13 AS=1.224e-13 PD=1.08e-06 PS=5.4e-07 w_cont=6e-07 nfing=1 mmm=1 $X=-197240 $Y=267620 $D=5
M51 gnd! vdd! gnd! cpoly_p w=3.8e-06 l=2e-06 c=5.2038e-14 as=2.31158e-13 ad=7.488e-13 ps=1.44e-06 pd=1.11673e-06 sim_w=2.88e-06 m_per_maxw=1.31944 numb_sub_cont=3 nfing=1 $X=-398620 $Y=276580 $D=21
M52 vdd! gnd! vdd! cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=-196800 $Y=283540 $D=22
M53 vdd! gnd! vdd! cpoly_n w=9.16e-06 l=2e-06 c=1.08961e-13 as=2.08643e-13 ad=1.4976e-12 ps=2.88e-06 pd=2.57123e-06 sim_w=5.76e-06 m_per_maxw=1.59028 numb_sub_cont=3 nfing=1 $X=-398400 $Y=283540 $D=22
R54 vdd! 21 454669 L=0.00067528 W=5e-07 m=1 $[rppoly] $X=-307340 $Y=260540 $D=19
R55 35 gnd! 636697 L=0.00094554 W=5e-07 m=1 $[rppoly] $X=-311920 $Y=-149700 $D=19
R56 gnd! 23 154847 L=0.00025532 W=5e-07 m=1 $[rppoly] $X=-432800 $Y=261340 $D=19
R57 58 41 618825 L=0.00091834 W=5e-07 m=1 $[rppoly] $X=-434020 $Y=-28040 $D=19
R58 41 vdd! 1.06273e+06 L=0.00157554 W=5e-07 m=1 $[rppoly] $X=-1013060 $Y=266360 $D=19
R59 15 47 198228 L=0.00029402 W=5e-07 m=1 $[rppoly] $X=-436800 $Y=265180 $D=19
R60 Usub 57 396298 L=0.00058782 W=5e-07 m=1 $[rppoly] $X=-435700 $Y=-28040 $D=19
R61 57 58 158908 L=0.00023598 W=5e-07 m=1 $[rppoly] $X=-434820 $Y=-147020 $D=19
D62 gnd! vdd! dn PJ=0.000409 m=1 $X=-395080 $Y=-149700 $D=8
D63 vdd! vdd! dn PJ=0.000409 m=1 $X=-392760 $Y=-149700 $D=8
D64 gnd! vdd! dn PJ=0.000409 m=1 $X=-385800 $Y=-149700 $D=8
D65 vdd! vdd! dn PJ=0.000409 m=1 $X=-383480 $Y=-149700 $D=8
D66 gnd! vdd! dn PJ=0.000409 m=1 $X=-376520 $Y=-149700 $D=8
D67 vdd! vdd! dn PJ=0.000409 m=1 $X=-374200 $Y=-149700 $D=8
D68 gnd! vdd! dn PJ=0.000409 m=1 $X=-367240 $Y=-149700 $D=8
D69 vdd! vdd! dn PJ=0.000409 m=1 $X=-364920 $Y=-149700 $D=8
D70 gnd! vdd! dn PJ=0.000409 m=1 $X=-357960 $Y=-149700 $D=8
D71 vdd! vdd! dn PJ=0.000409 m=1 $X=-355640 $Y=-149700 $D=8
D72 gnd! vdd! dn PJ=0.000409 m=1 $X=-348680 $Y=-149700 $D=8
D73 vdd! vdd! dn PJ=0.000409 m=1 $X=-346360 $Y=-149700 $D=8
D74 gnd! vdd! dn PJ=0.000409 m=1 $X=-339400 $Y=-149700 $D=8
D75 vdd! vdd! dn PJ=0.000409 m=1 $X=-337080 $Y=-149700 $D=8
D76 gnd! vdd! dn PJ=0.000409 m=1 $X=-330120 $Y=-149700 $D=8
D77 vdd! vdd! dn PJ=0.000409 m=1 $X=-327800 $Y=-149700 $D=8
D78 gnd! vdd! dn PJ=0.000409 m=1 $X=-320840 $Y=-149700 $D=8
D79 vdd! vdd! dn PJ=0.000409 m=1 $X=-318520 $Y=-149700 $D=8
D80 gnd! vdd! dn PJ=0.000409 m=1 $X=-432200 $Y=-149700 $D=8
D81 vdd! vdd! dn PJ=0.000409 m=1 $X=-429880 $Y=-149700 $D=8
D82 gnd! vdd! dn PJ=0.000409 m=1 $X=-422920 $Y=-149700 $D=8
D83 vdd! vdd! dn PJ=0.000409 m=1 $X=-420600 $Y=-149700 $D=8
D84 gnd! vdd! dn PJ=0.000409 m=1 $X=-413640 $Y=-149700 $D=8
D85 vdd! vdd! dn PJ=0.000409 m=1 $X=-411320 $Y=-149700 $D=8
D86 gnd! vdd! dn PJ=0.000409 m=1 $X=-404360 $Y=-149700 $D=8
D87 vdd! vdd! dn PJ=0.000409 m=1 $X=-402040 $Y=-149700 $D=8
D88 gnd! vdd! dn PJ=0.000409 m=1 $X=-398100 $Y=-149700 $D=9
D89 vdd! vdd! dn PJ=0.000409 m=1 $X=-391140 $Y=-149700 $D=9
D90 gnd! vdd! dn PJ=0.000409 m=1 $X=-388820 $Y=-149700 $D=9
D91 vdd! vdd! dn PJ=0.000409 m=1 $X=-381860 $Y=-149700 $D=9
D92 gnd! vdd! dn PJ=0.000409 m=1 $X=-379540 $Y=-149700 $D=9
D93 vdd! vdd! dn PJ=0.000409 m=1 $X=-372580 $Y=-149700 $D=9
D94 gnd! vdd! dn PJ=0.000409 m=1 $X=-370260 $Y=-149700 $D=9
D95 vdd! vdd! dn PJ=0.000409 m=1 $X=-363300 $Y=-149700 $D=9
D96 gnd! vdd! dn PJ=0.000409 m=1 $X=-360980 $Y=-149700 $D=9
D97 vdd! vdd! dn PJ=0.000409 m=1 $X=-354020 $Y=-149700 $D=9
D98 gnd! vdd! dn PJ=0.000409 m=1 $X=-351700 $Y=-149700 $D=9
D99 vdd! vdd! dn PJ=0.000409 m=1 $X=-344740 $Y=-149700 $D=9
D100 gnd! vdd! dn PJ=0.000409 m=1 $X=-342420 $Y=-149700 $D=9
D101 vdd! vdd! dn PJ=0.000409 m=1 $X=-335460 $Y=-149700 $D=9
D102 gnd! vdd! dn PJ=0.000409 m=1 $X=-333140 $Y=-149700 $D=9
D103 vdd! vdd! dn PJ=0.000409 m=1 $X=-326180 $Y=-149700 $D=9
D104 gnd! vdd! dn PJ=0.000409 m=1 $X=-323860 $Y=-149700 $D=9
D105 vdd! vdd! dn PJ=0.000409 m=1 $X=-316900 $Y=-149700 $D=9
D106 gnd! vdd! dn PJ=0.000409 m=1 $X=-314580 $Y=-149700 $D=9
D107 vdd! vdd! dn PJ=0.000409 m=1 $X=-428260 $Y=-149700 $D=9
D108 gnd! vdd! dn PJ=0.000409 m=1 $X=-425940 $Y=-149700 $D=9
D109 vdd! vdd! dn PJ=0.000409 m=1 $X=-418980 $Y=-149700 $D=9
D110 gnd! vdd! dn PJ=0.000409 m=1 $X=-416660 $Y=-149700 $D=9
D111 vdd! vdd! dn PJ=0.000409 m=1 $X=-409700 $Y=-149700 $D=9
D112 gnd! vdd! dn PJ=0.000409 m=1 $X=-407380 $Y=-149700 $D=9
D113 vdd! vdd! dn PJ=0.000409 m=1 $X=-400420 $Y=-149700 $D=9
X114 gnd! Usub 14 15 17 18 19 ICV_94 $T=-437300 -146840 1 180 $X=-451980 $Y=-150000
X115 gnd! Usub 14 15 17 18 19 ICV_95 $T=-451980 -146840 1 180 $X=-466660 $Y=-150000
X116 gnd! Usub 14 15 17 18 19 ICV_96 $T=-466660 -146840 1 180 $X=-481340 $Y=-150000
X117 gnd! Usub 14 15 17 18 19 ICV_97 $T=-481340 -146840 1 180 $X=-496020 $Y=-150000
X118 gnd! Usub 14 15 17 18 19 ICV_98 $T=-496020 -146840 1 180 $X=-510700 $Y=-150000
X119 gnd! Usub 14 15 17 18 19 ICV_99 $T=-510700 -146840 1 180 $X=-525380 $Y=-150000
X120 gnd! Usub 14 15 17 18 19 ICV_100 $T=-525380 -146840 1 180 $X=-540060 $Y=-150000
X121 gnd! Usub 14 15 17 18 19 ICV_101 $T=-540060 -146840 1 180 $X=-554740 $Y=-150000
X122 gnd! Usub 14 15 17 18 19 ICV_102 $T=-554740 -146840 1 180 $X=-569420 $Y=-150000
X123 gnd! Usub 14 15 17 18 19 ICV_103 $T=-569420 -146840 1 180 $X=-584100 $Y=-150000
X124 gnd! Usub 14 15 17 18 19 ICV_104 $T=-584100 -146840 1 180 $X=-598780 $Y=-150000
X125 gnd! Usub 14 15 17 18 19 ICV_105 $T=-598780 -146840 1 180 $X=-613460 $Y=-150000
X126 gnd! Usub 14 15 17 18 19 ICV_106 $T=-613460 -146840 1 180 $X=-628140 $Y=-150000
X127 gnd! Usub 14 15 17 18 19 ICV_107 $T=-628140 -146840 1 180 $X=-642820 $Y=-150000
X128 gnd! Usub 14 15 17 18 19 ICV_108 $T=-642820 -146840 1 180 $X=-657500 $Y=-150000
X129 gnd! Usub 14 15 17 18 19 ICV_109 $T=-657500 -146840 1 180 $X=-672180 $Y=-150000
X130 gnd! Usub 14 15 17 18 19 ICV_110 $T=-672180 -146840 1 180 $X=-686860 $Y=-150000
X131 gnd! Usub 14 15 17 18 19 ICV_111 $T=-686860 -146840 1 180 $X=-701540 $Y=-150000
X132 gnd! Usub 14 15 17 18 19 ICV_112 $T=-701540 -146840 1 180 $X=-716220 $Y=-150000
X133 gnd! Usub 14 15 17 18 19 ICV_113 $T=-716220 -146840 1 180 $X=-730900 $Y=-150000
X134 gnd! Usub 14 15 17 18 19 ICV_114 $T=-730900 -146840 1 180 $X=-745580 $Y=-150000
X135 gnd! Usub 14 15 17 18 19 ICV_115 $T=-745580 -146840 1 180 $X=-760260 $Y=-150000
X136 gnd! Usub 14 15 17 18 19 ICV_116 $T=-760260 -146840 1 180 $X=-774940 $Y=-150000
X137 gnd! Usub 14 15 17 18 19 ICV_117 $T=-774940 -146840 1 180 $X=-789620 $Y=-150000
X138 gnd! Usub 14 15 17 18 19 ICV_118 $T=-789620 -146840 1 180 $X=-804300 $Y=-150000
X139 gnd! Usub 14 15 17 18 19 ICV_119 $T=-804300 -146840 1 180 $X=-818980 $Y=-150000
X140 gnd! Usub 14 15 17 18 19 ICV_120 $T=-818980 -146840 1 180 $X=-833660 $Y=-150000
X141 gnd! Usub 14 15 17 18 19 ICV_121 $T=-833660 -146840 1 180 $X=-848340 $Y=-150000
X142 gnd! Usub 14 15 17 18 19 ICV_122 $T=-848340 -146840 1 180 $X=-863020 $Y=-150000
X143 gnd! Usub 14 15 17 18 19 ICV_123 $T=-863020 -146840 1 180 $X=-877700 $Y=-150000
X144 gnd! Usub 14 15 17 18 19 ICV_124 $T=-877700 -146840 1 180 $X=-892380 $Y=-150000
X145 gnd! Usub 14 15 17 18 19 ICV_125 $T=-892380 -146840 1 180 $X=-907060 $Y=-150000
X146 gnd! Usub 14 15 17 18 19 ICV_126 $T=-907060 -146840 1 180 $X=-921740 $Y=-150000
X147 gnd! Usub 14 15 17 18 19 ICV_127 $T=-921740 -146840 1 180 $X=-936420 $Y=-150000
X148 gnd! Usub 14 15 17 18 19 ICV_128 $T=-936420 -146840 1 180 $X=-951100 $Y=-150000
X149 gnd! Usub 14 15 17 18 19 ICV_129 $T=-951100 -146840 1 180 $X=-965780 $Y=-150000
X150 gnd! Usub 14 15 17 18 19 ICV_130 $T=-965780 -146840 1 180 $X=-980460 $Y=-150000
X151 gnd! Usub 14 15 17 18 19 ICV_131 $T=-980460 -146840 1 180 $X=-995140 $Y=-150000
X152 gnd! Usub 14 15 17 18 19 ICV_132 $T=-995140 -146840 1 180 $X=-1009820 $Y=-150000
X153 gnd! vdd! 20 21 26 25 24 27 30 53 28 29 ICV_133 $T=0 0 0 0 $X=-195500 $Y=268500
X154 gnd! vdd! 30 49 28 29 33 ICV_136 $T=0 0 0 0 $X=-195500 $Y=159400
X155 30 33 ICV_139 $T=0 0 0 0 $X=-195500 $Y=61280
X156 gnd! 15 17 31 33 32 54 14 55 34 ICV_144 $T=0 0 0 0 $X=-195500 $Y=-37700
X157 14 36 ICV_147 $T=0 0 0 0 $X=-195500 $Y=-143200
X158 17 36 14 35 ICV_148 $T=0 0 0 0 $X=-195500 $Y=-286000
X159 gnd! vdd! 23 21 20 24 40 39 41 42 43 44 22 56 45 25 38 37 ICV_151 $T=0 0 0 0 $X=-398300 $Y=268020
X160 gnd! vdd! 23 20 22 41 40 42 43 44 51 34 ICV_152 $T=0 0 0 0 $X=-398300 $Y=159400
X161 22 34 ICV_153 $T=0 0 0 0 $X=-398300 $Y=61280
X162 gnd! 17 15 54 55 14 34 31 32 33 ICV_154 $T=0 0 0 0 $X=-398300 $Y=-37700
X163 14 36 ICV_155 $T=0 0 0 0 $X=-398300 $Y=-143200
X164 17 36 35 14 ICV_156 $T=0 0 0 0 $X=-398300 $Y=-286000
X165 nTest gnd! vdd! 46 38 39 37 40 ICV_160 $T=0 0 0 0 $X=-1015000 $Y=268500
X168 Usub 47 14 ICV_163 $T=0 0 0 0 $X=-1015000 $Y=-37700
X169 Usub 14 48 47 ICV_164 $T=0 0 0 0 $X=-1015000 $Y=-146960
.ENDS
***************************************
.SUBCKT ICV_166 1 2
** N=5 EP=2 IP=8 FDC=3576
X0 1 2 Fill_Block_8Kx8 $T=-440480 0 0 0 $X=-440840 $Y=-320
X1 1 2 Fill_Block_8Kx8 $T=0 0 0 0 $X=-360 $Y=-320
.ENDS
***************************************
.SUBCKT ICV_167 1 2
** N=5 EP=2 IP=8 FDC=7152
X0 1 2 ICV_166 $T=-880960 0 0 0 $X=-1321800 $Y=-320
X1 1 2 ICV_166 $T=0 0 0 0 $X=-440840 $Y=-320
.ENDS
***************************************
.SUBCKT RingPad DO_Bank<1> DI_Bank<1> DO_Bank<2> DI_Bank<2> DO_Bank<3> DI_Bank<3> DO_Bank<4> DI_Bank<4> DO_Bank<5> Adr<0> DI_Bank<5> DO_Bank<7> Adr<1> DO_Bank<6> DI_Bank<6> Adr<2> Adr<3> DI_Bank<7> DO_Bank<8> DI_Bank<8>
+ Adr<4> DO_Bank<17> Adr<5> DI_Bank<17> Adr<6> DO_Bank<18> Adr<7> DI_Bank<18> DO_Bank<19> DI_Bank<19> DO_Bank<20> DI_Bank<20> DO_Bank<21> DI_Bank<21> Adr<8> DO_Bank<23> Adr<9> DO_Bank<22> DI_Bank<22> Adr<10>
+ DI_Bank<23> DO_Bank<24> DI_Bank<24> Bit_16 Bit_32 nCE nOE_Core nWE Adr<12> Adr<19> Adr<18> Adr<17> DI_Bank<9> Adr<11> DI_Bank<10> DO_Bank<9> DI_Bank<11> DO_Bank<10> DO_Bank<11> DI_Bank<12>
+ DO_Bank<12> DI_Bank<13> DO_Bank<13> DI_Bank<14> DO_Bank<14> DI_Bank<15> DO_Bank<15> DI_Bank<16> Adr<13> DO_Bank<16> Adr<14> DI_Bank<25> Adr<15> DI_Bank<26> DO_Bank<25> Adr<16> DI_Bank<27> DO_Bank<26> DI_Bank<28> DO_Bank<27>
+ DO_Bank<28> DI_Bank<29> DO_Bank<29> DI_Bank<30> DO_Bank<30> DI_Bank<31> DO_Bank<31> DI_Bank<32> DO_Bank<32> GND_PAD! VDD_PAD! gnd! vdd! NWR BIT32 BIT16 DIO5 DIO21 DIO13 DIO29
+ DIO8 DIO24 DIO16 DIO32 DIO2 DIO1 DIO4 DIO3 DIO7 DIO6 DIO18 DIO17 DIO20 DIO19 DIO23 DIO22 DIO10 DIO9 DIO12 DIO11
+ DIO15 DIO14 DIO26 DIO25 DIO28 DIO27 DIO31 DIO30 A18 A19 A0 A1 A2 A3 A4 A5 A6 A7 A8 A9
+ A10 A11 A12 A13 A14 A15 A16 A17 OEN CEN Test MODE A20 CS1 CS2 A21 Usub
** N=698 EP=157 IP=1830 FDC=351497
M0 1 534 gnd! gnd! nmos_a L=2.4e-07 W=2.4e-06 AD=1.4e-12 AS=9.6e-13 PD=3.5e-06 PS=1.75e-06 w_cont=1.1e-06 nfing=1 source_num=2 $X=11640 $Y=13210580 $D=1
M1 154 584 gnd! gnd! nmos_a L=2.4e-07 W=2.4e-06 AD=1.4e-12 AS=9.6e-13 PD=3.5e-06 PS=1.75e-06 w_cont=1.1e-06 nfing=1 source_num=2 $X=14079000 $Y=13210580 $D=1
M2 97 98 gnd! gnd! nmos_a L=2.4e-07 W=1.2e-06 AD=4.68e-13 AS=4.8e-13 PD=9e-07 PS=9e-07 w_cont=6e-07 nfing=1 source_num=2 $X=7799080 $Y=13213660 $D=1
M3 97 563 gnd! gnd! nmos_a L=2.4e-07 W=1.2e-06 AD=4.68e-13 AS=4.8e-13 PD=9e-07 PS=9e-07 w_cont=6e-07 nfing=1 source_num=2 $X=7799840 $Y=13213660 $D=1
M4 97 98 562 562 pmos_a L=2.4e-07 W=2.4e-06 AD=1.2e-12 AS=1.32e-13 PD=3e-06 PS=1.5e-06 w_cont=6e-07 nfing=1 mmm=1 $X=7799080 $Y=13208060 $D=5
M5 562 563 vdd! vdd! pmos_a L=2.4e-07 W=2.4e-06 AD=1.2e-12 AS=1.68e-13 PD=3e-06 PS=1.5e-06 w_cont=6e-07 nfing=1 mmm=1 $X=7800520 $Y=13208060 $D=5
M6 98 697 vdd! vdd! pmos_a L=2.4e-07 W=2.4e-06 AD=7.8e-13 AS=1.32e-13 PD=1.5e-06 PS=1.5e-06 w_cont=6e-07 nfing=1 mmm=1 $X=6558480 $Y=13208060 $D=5
M7 563 698 vdd! vdd! pmos_a L=2.4e-07 W=2.4e-06 AD=7.8e-13 AS=1.68e-13 PD=1.5e-06 PS=1.5e-06 w_cont=6e-07 nfing=1 mmm=1 $X=7801280 $Y=13208060 $D=5
D8 GND_PAD! VDD_PAD! dn PJ=0.00041 m=1 $X=-38460 $Y=80300 $D=8
D9 GND_PAD! VDD_PAD! dn PJ=0.00041 m=1 $X=-28460 $Y=80300 $D=8
D10 GND_PAD! VDD_PAD! dn PJ=0.00041 m=1 $X=-18460 $Y=80300 $D=8
D11 GND_PAD! VDD_PAD! dn PJ=0.00041 m=1 $X=-8460 $Y=80300 $D=8
D12 GND_PAD! VDD_PAD! dn PJ=0.00041 m=1 $X=1540 $Y=80300 $D=8
D13 GND_PAD! VDD_PAD! dn PJ=0.00041 m=1 $X=11540 $Y=80300 $D=8
D14 GND_PAD! VDD_PAD! dn PJ=0.00041 m=1 $X=21540 $Y=80300 $D=8
D15 GND_PAD! VDD_PAD! dn PJ=0.00041 m=1 $X=31540 $Y=80300 $D=8
D16 GND_PAD! VDD_PAD! dn PJ=0.00041 m=1 $X=41540 $Y=80300 $D=8
D17 MODE vdd! dn PJ=0.0002 m=1 $X=1024020 $Y=13228100 $D=8
D18 MODE vdd! dn PJ=0.0002 m=1 $X=1024020 $Y=13438100 $D=8
D19 gnd! MODE dn PJ=0.0002 m=1 $X=1026340 $Y=13232500 $D=8
D20 gnd! MODE dn PJ=0.0002 m=1 $X=1026340 $Y=13442500 $D=8
D21 MODE vdd! dn PJ=0.0002 m=1 $X=1028660 $Y=13228100 $D=8
D22 MODE vdd! dn PJ=0.0002 m=1 $X=1028660 $Y=13438100 $D=8
D23 gnd! MODE dn PJ=0.0001 m=1 $X=1030980 $Y=13332500 $D=8
D24 gnd! MODE dn PJ=0.0001 m=1 $X=1030980 $Y=13542500 $D=8
D25 MODE vdd! dn PJ=0.0001 m=1 $X=1034160 $Y=13228100 $D=8
D26 MODE vdd! dn PJ=0.0001 m=1 $X=1034160 $Y=13438100 $D=8
D27 gnd! MODE dn PJ=0.0002 m=1 $X=1036480 $Y=13232500 $D=8
D28 gnd! MODE dn PJ=0.0002 m=1 $X=1036480 $Y=13442500 $D=8
D29 MODE vdd! dn PJ=0.0002 m=1 $X=1038800 $Y=13228100 $D=8
D30 MODE vdd! dn PJ=0.0002 m=1 $X=1038800 $Y=13438100 $D=8
D31 gnd! MODE dn PJ=0.0002 m=1 $X=1041120 $Y=13232500 $D=8
D32 gnd! MODE dn PJ=0.0002 m=1 $X=1041120 $Y=13442500 $D=8
D33 MODE vdd! dn PJ=0.0002 m=1 $X=1043440 $Y=13228100 $D=8
D34 MODE vdd! dn PJ=0.0002 m=1 $X=1043440 $Y=13438100 $D=8
D35 gnd! MODE dn PJ=0.0001 m=1 $X=1045760 $Y=13332500 $D=8
D36 gnd! MODE dn PJ=0.0001 m=1 $X=1045760 $Y=13542500 $D=8
D37 MODE vdd! dn PJ=0.0001 m=1 $X=1048940 $Y=13228100 $D=8
D38 MODE vdd! dn PJ=0.0001 m=1 $X=1048940 $Y=13438100 $D=8
D39 gnd! MODE dn PJ=0.0002 m=1 $X=1051260 $Y=13232500 $D=8
D40 gnd! MODE dn PJ=0.0002 m=1 $X=1051260 $Y=13442500 $D=8
D41 MODE vdd! dn PJ=0.0002 m=1 $X=1053580 $Y=13228100 $D=8
D42 MODE vdd! dn PJ=0.0002 m=1 $X=1053580 $Y=13438100 $D=8
D43 gnd! MODE dn PJ=0.0002 m=1 $X=1055900 $Y=13232500 $D=8
D44 gnd! MODE dn PJ=0.0002 m=1 $X=1055900 $Y=13442500 $D=8
D45 MODE vdd! dn PJ=0.0002 m=1 $X=1058220 $Y=13228100 $D=8
D46 MODE vdd! dn PJ=0.0002 m=1 $X=1058220 $Y=13438100 $D=8
D47 gnd! MODE dn PJ=0.0001 m=1 $X=1060540 $Y=13332500 $D=8
D48 gnd! MODE dn PJ=0.0001 m=1 $X=1060540 $Y=13542500 $D=8
D49 MODE vdd! dn PJ=0.0001 m=1 $X=1063720 $Y=13228100 $D=8
D50 MODE vdd! dn PJ=0.0001 m=1 $X=1063720 $Y=13438100 $D=8
D51 gnd! MODE dn PJ=0.0002 m=1 $X=1066040 $Y=13232500 $D=8
D52 gnd! MODE dn PJ=0.0002 m=1 $X=1066040 $Y=13442500 $D=8
D53 MODE vdd! dn PJ=0.0002 m=1 $X=1068360 $Y=13228100 $D=8
D54 MODE vdd! dn PJ=0.0002 m=1 $X=1068360 $Y=13438100 $D=8
D55 gnd! MODE dn PJ=0.0002 m=1 $X=1070680 $Y=13232500 $D=8
D56 gnd! MODE dn PJ=0.0002 m=1 $X=1070680 $Y=13442500 $D=8
D57 MODE vdd! dn PJ=0.0002 m=1 $X=1073000 $Y=13228100 $D=8
D58 MODE vdd! dn PJ=0.0002 m=1 $X=1073000 $Y=13438100 $D=8
D59 gnd! MODE dn PJ=0.0001 m=1 $X=1075320 $Y=13332500 $D=8
D60 gnd! MODE dn PJ=0.0001 m=1 $X=1075320 $Y=13542500 $D=8
D61 MODE vdd! dn PJ=0.0001 m=1 $X=1078500 $Y=13228100 $D=8
D62 MODE vdd! dn PJ=0.0001 m=1 $X=1078500 $Y=13438100 $D=8
D63 gnd! MODE dn PJ=0.0002 m=1 $X=1080820 $Y=13232500 $D=8
D64 gnd! MODE dn PJ=0.0002 m=1 $X=1080820 $Y=13442500 $D=8
D65 MODE vdd! dn PJ=0.0002 m=1 $X=1083140 $Y=13228100 $D=8
D66 MODE vdd! dn PJ=0.0002 m=1 $X=1083140 $Y=13438100 $D=8
D67 gnd! MODE dn PJ=0.0002 m=1 $X=1085460 $Y=13232500 $D=8
D68 gnd! MODE dn PJ=0.0002 m=1 $X=1085460 $Y=13442500 $D=8
D69 MODE vdd! dn PJ=0.0002 m=1 $X=1087780 $Y=13228100 $D=8
D70 MODE vdd! dn PJ=0.0002 m=1 $X=1087780 $Y=13438100 $D=8
D71 gnd! MODE dn PJ=0.0001 m=1 $X=1090100 $Y=13332500 $D=8
D72 gnd! MODE dn PJ=0.0001 m=1 $X=1090100 $Y=13542500 $D=8
D73 MODE vdd! dn PJ=0.0001 m=1 $X=1093280 $Y=13228100 $D=8
D74 MODE vdd! dn PJ=0.0001 m=1 $X=1093280 $Y=13438100 $D=8
D75 gnd! MODE dn PJ=0.0002 m=1 $X=1095600 $Y=13232500 $D=8
D76 gnd! MODE dn PJ=0.0002 m=1 $X=1095600 $Y=13442500 $D=8
D77 MODE vdd! dn PJ=0.0002 m=1 $X=1097920 $Y=13228100 $D=8
D78 MODE vdd! dn PJ=0.0002 m=1 $X=1097920 $Y=13438100 $D=8
D79 gnd! MODE dn PJ=0.0002 m=1 $X=1100240 $Y=13232500 $D=8
D80 gnd! MODE dn PJ=0.0002 m=1 $X=1100240 $Y=13442500 $D=8
D81 MODE vdd! dn PJ=0.0002 m=1 $X=1102560 $Y=13228100 $D=8
D82 MODE vdd! dn PJ=0.0002 m=1 $X=1102560 $Y=13438100 $D=8
D83 gnd! MODE dn PJ=0.0001 m=1 $X=1104880 $Y=13332500 $D=8
D84 gnd! MODE dn PJ=0.0001 m=1 $X=1104880 $Y=13542500 $D=8
D85 MODE vdd! dn PJ=0.0001 m=1 $X=1108060 $Y=13228100 $D=8
D86 MODE vdd! dn PJ=0.0001 m=1 $X=1108060 $Y=13438100 $D=8
D87 gnd! MODE dn PJ=0.0002 m=1 $X=1110380 $Y=13232500 $D=8
D88 gnd! MODE dn PJ=0.0002 m=1 $X=1110380 $Y=13442500 $D=8
D89 MODE vdd! dn PJ=0.0002 m=1 $X=1112700 $Y=13228100 $D=8
D90 MODE vdd! dn PJ=0.0002 m=1 $X=1112700 $Y=13438100 $D=8
D91 gnd! MODE dn PJ=0.0002 m=1 $X=1115020 $Y=13232500 $D=8
D92 gnd! MODE dn PJ=0.0002 m=1 $X=1115020 $Y=13442500 $D=8
D93 A2 vdd! dn PJ=0.0002 m=1 $X=2324020 $Y=13228100 $D=8
D94 A2 vdd! dn PJ=0.0002 m=1 $X=2324020 $Y=13438100 $D=8
D95 gnd! A2 dn PJ=0.0002 m=1 $X=2326340 $Y=13232500 $D=8
D96 gnd! A2 dn PJ=0.0002 m=1 $X=2326340 $Y=13442500 $D=8
D97 A2 vdd! dn PJ=0.0002 m=1 $X=2328660 $Y=13228100 $D=8
D98 A2 vdd! dn PJ=0.0002 m=1 $X=2328660 $Y=13438100 $D=8
D99 gnd! A2 dn PJ=0.0001 m=1 $X=2330980 $Y=13332500 $D=8
D100 gnd! A2 dn PJ=0.0001 m=1 $X=2330980 $Y=13542500 $D=8
D101 A2 vdd! dn PJ=0.0001 m=1 $X=2334160 $Y=13228100 $D=8
D102 A2 vdd! dn PJ=0.0001 m=1 $X=2334160 $Y=13438100 $D=8
D103 gnd! A2 dn PJ=0.0002 m=1 $X=2336480 $Y=13232500 $D=8
D104 gnd! A2 dn PJ=0.0002 m=1 $X=2336480 $Y=13442500 $D=8
D105 A2 vdd! dn PJ=0.0002 m=1 $X=2338800 $Y=13228100 $D=8
D106 A2 vdd! dn PJ=0.0002 m=1 $X=2338800 $Y=13438100 $D=8
D107 gnd! A2 dn PJ=0.0002 m=1 $X=2341120 $Y=13232500 $D=8
D108 gnd! A2 dn PJ=0.0002 m=1 $X=2341120 $Y=13442500 $D=8
D109 A2 vdd! dn PJ=0.0002 m=1 $X=2343440 $Y=13228100 $D=8
D110 A2 vdd! dn PJ=0.0002 m=1 $X=2343440 $Y=13438100 $D=8
D111 gnd! A2 dn PJ=0.0001 m=1 $X=2345760 $Y=13332500 $D=8
D112 gnd! A2 dn PJ=0.0001 m=1 $X=2345760 $Y=13542500 $D=8
D113 A2 vdd! dn PJ=0.0001 m=1 $X=2348940 $Y=13228100 $D=8
D114 A2 vdd! dn PJ=0.0001 m=1 $X=2348940 $Y=13438100 $D=8
D115 gnd! A2 dn PJ=0.0002 m=1 $X=2351260 $Y=13232500 $D=8
D116 gnd! A2 dn PJ=0.0002 m=1 $X=2351260 $Y=13442500 $D=8
D117 A2 vdd! dn PJ=0.0002 m=1 $X=2353580 $Y=13228100 $D=8
D118 A2 vdd! dn PJ=0.0002 m=1 $X=2353580 $Y=13438100 $D=8
D119 gnd! A2 dn PJ=0.0002 m=1 $X=2355900 $Y=13232500 $D=8
D120 gnd! A2 dn PJ=0.0002 m=1 $X=2355900 $Y=13442500 $D=8
D121 A2 vdd! dn PJ=0.0002 m=1 $X=2358220 $Y=13228100 $D=8
D122 A2 vdd! dn PJ=0.0002 m=1 $X=2358220 $Y=13438100 $D=8
D123 gnd! A2 dn PJ=0.0001 m=1 $X=2360540 $Y=13332500 $D=8
D124 gnd! A2 dn PJ=0.0001 m=1 $X=2360540 $Y=13542500 $D=8
D125 A2 vdd! dn PJ=0.0001 m=1 $X=2363720 $Y=13228100 $D=8
D126 A2 vdd! dn PJ=0.0001 m=1 $X=2363720 $Y=13438100 $D=8
D127 gnd! A2 dn PJ=0.0002 m=1 $X=2366040 $Y=13232500 $D=8
D128 gnd! A2 dn PJ=0.0002 m=1 $X=2366040 $Y=13442500 $D=8
D129 A2 vdd! dn PJ=0.0002 m=1 $X=2368360 $Y=13228100 $D=8
D130 A2 vdd! dn PJ=0.0002 m=1 $X=2368360 $Y=13438100 $D=8
D131 gnd! A2 dn PJ=0.0002 m=1 $X=2370680 $Y=13232500 $D=8
D132 gnd! A2 dn PJ=0.0002 m=1 $X=2370680 $Y=13442500 $D=8
D133 A2 vdd! dn PJ=0.0002 m=1 $X=2373000 $Y=13228100 $D=8
D134 A2 vdd! dn PJ=0.0002 m=1 $X=2373000 $Y=13438100 $D=8
D135 gnd! A2 dn PJ=0.0001 m=1 $X=2375320 $Y=13332500 $D=8
D136 gnd! A2 dn PJ=0.0001 m=1 $X=2375320 $Y=13542500 $D=8
D137 A2 vdd! dn PJ=0.0001 m=1 $X=2378500 $Y=13228100 $D=8
D138 A2 vdd! dn PJ=0.0001 m=1 $X=2378500 $Y=13438100 $D=8
D139 gnd! A2 dn PJ=0.0002 m=1 $X=2380820 $Y=13232500 $D=8
D140 gnd! A2 dn PJ=0.0002 m=1 $X=2380820 $Y=13442500 $D=8
D141 A2 vdd! dn PJ=0.0002 m=1 $X=2383140 $Y=13228100 $D=8
D142 A2 vdd! dn PJ=0.0002 m=1 $X=2383140 $Y=13438100 $D=8
D143 gnd! A2 dn PJ=0.0002 m=1 $X=2385460 $Y=13232500 $D=8
D144 gnd! A2 dn PJ=0.0002 m=1 $X=2385460 $Y=13442500 $D=8
D145 A2 vdd! dn PJ=0.0002 m=1 $X=2387780 $Y=13228100 $D=8
D146 A2 vdd! dn PJ=0.0002 m=1 $X=2387780 $Y=13438100 $D=8
D147 gnd! A2 dn PJ=0.0001 m=1 $X=2390100 $Y=13332500 $D=8
D148 gnd! A2 dn PJ=0.0001 m=1 $X=2390100 $Y=13542500 $D=8
D149 A2 vdd! dn PJ=0.0001 m=1 $X=2393280 $Y=13228100 $D=8
D150 A2 vdd! dn PJ=0.0001 m=1 $X=2393280 $Y=13438100 $D=8
D151 gnd! A2 dn PJ=0.0002 m=1 $X=2395600 $Y=13232500 $D=8
D152 gnd! A2 dn PJ=0.0002 m=1 $X=2395600 $Y=13442500 $D=8
D153 A2 vdd! dn PJ=0.0002 m=1 $X=2397920 $Y=13228100 $D=8
D154 A2 vdd! dn PJ=0.0002 m=1 $X=2397920 $Y=13438100 $D=8
D155 gnd! A2 dn PJ=0.0002 m=1 $X=2400240 $Y=13232500 $D=8
D156 gnd! A2 dn PJ=0.0002 m=1 $X=2400240 $Y=13442500 $D=8
D157 A2 vdd! dn PJ=0.0002 m=1 $X=2402560 $Y=13228100 $D=8
D158 A2 vdd! dn PJ=0.0002 m=1 $X=2402560 $Y=13438100 $D=8
D159 gnd! A2 dn PJ=0.0001 m=1 $X=2404880 $Y=13332500 $D=8
D160 gnd! A2 dn PJ=0.0001 m=1 $X=2404880 $Y=13542500 $D=8
D161 A2 vdd! dn PJ=0.0001 m=1 $X=2408060 $Y=13228100 $D=8
D162 A2 vdd! dn PJ=0.0001 m=1 $X=2408060 $Y=13438100 $D=8
D163 gnd! A2 dn PJ=0.0002 m=1 $X=2410380 $Y=13232500 $D=8
D164 gnd! A2 dn PJ=0.0002 m=1 $X=2410380 $Y=13442500 $D=8
D165 A2 vdd! dn PJ=0.0002 m=1 $X=2412700 $Y=13228100 $D=8
D166 A2 vdd! dn PJ=0.0002 m=1 $X=2412700 $Y=13438100 $D=8
D167 gnd! A2 dn PJ=0.0002 m=1 $X=2415020 $Y=13232500 $D=8
D168 gnd! A2 dn PJ=0.0002 m=1 $X=2415020 $Y=13442500 $D=8
D169 GND_PAD! VDD_PAD! dn PJ=0.00041 m=1 $X=3261540 $Y=80300 $D=8
D170 GND_PAD! VDD_PAD! dn PJ=0.00041 m=1 $X=3271540 $Y=80300 $D=8
D171 GND_PAD! VDD_PAD! dn PJ=0.00041 m=1 $X=3281540 $Y=80300 $D=8
D172 GND_PAD! VDD_PAD! dn PJ=0.00041 m=1 $X=3291540 $Y=80300 $D=8
D173 GND_PAD! VDD_PAD! dn PJ=0.00041 m=1 $X=3301540 $Y=80300 $D=8
D174 GND_PAD! VDD_PAD! dn PJ=0.00041 m=1 $X=3311540 $Y=80300 $D=8
D175 GND_PAD! VDD_PAD! dn PJ=0.00041 m=1 $X=3321540 $Y=80300 $D=8
D176 GND_PAD! VDD_PAD! dn PJ=0.00041 m=1 $X=3331540 $Y=80300 $D=8
D177 GND_PAD! VDD_PAD! dn PJ=0.00041 m=1 $X=3341540 $Y=80300 $D=8
D178 VDD_PAD! vdd! dn PJ=0.00041 m=1 $X=3551760 $Y=80300 $D=8
D179 GND_PAD! VDD_PAD! dn PJ=0.00041 m=1 $X=3554260 $Y=80300 $D=8
D180 vdd! VDD_PAD! dn PJ=0.00041 m=1 $X=3559260 $Y=80300 $D=8
D181 VDD_PAD! vdd! dn PJ=0.00041 m=1 $X=3561760 $Y=80300 $D=8
D182 GND_PAD! VDD_PAD! dn PJ=0.00041 m=1 $X=3564260 $Y=80300 $D=8
D183 vdd! VDD_PAD! dn PJ=0.00041 m=1 $X=3569260 $Y=80300 $D=8
D184 VDD_PAD! vdd! dn PJ=0.00041 m=1 $X=3571760 $Y=80300 $D=8
D185 GND_PAD! VDD_PAD! dn PJ=0.00041 m=1 $X=3574260 $Y=80300 $D=8
D186 vdd! VDD_PAD! dn PJ=0.00041 m=1 $X=3579260 $Y=80300 $D=8
D187 VDD_PAD! vdd! dn PJ=0.00041 m=1 $X=3581760 $Y=80300 $D=8
D188 GND_PAD! VDD_PAD! dn PJ=0.00041 m=1 $X=3584260 $Y=80300 $D=8
D189 vdd! VDD_PAD! dn PJ=0.00041 m=1 $X=3589260 $Y=80300 $D=8
D190 VDD_PAD! vdd! dn PJ=0.00041 m=1 $X=3591760 $Y=80300 $D=8
D191 GND_PAD! VDD_PAD! dn PJ=0.00041 m=1 $X=3594260 $Y=80300 $D=8
D192 vdd! VDD_PAD! dn PJ=0.00041 m=1 $X=3599260 $Y=80300 $D=8
D193 VDD_PAD! vdd! dn PJ=0.00041 m=1 $X=3601760 $Y=80300 $D=8
D194 GND_PAD! VDD_PAD! dn PJ=0.00041 m=1 $X=3604260 $Y=80300 $D=8
D195 vdd! VDD_PAD! dn PJ=0.00041 m=1 $X=3609260 $Y=80300 $D=8
D196 VDD_PAD! vdd! dn PJ=0.00041 m=1 $X=3611760 $Y=80300 $D=8
D197 GND_PAD! VDD_PAD! dn PJ=0.00041 m=1 $X=3614260 $Y=80300 $D=8
D198 vdd! VDD_PAD! dn PJ=0.00041 m=1 $X=3619260 $Y=80300 $D=8
D199 VDD_PAD! vdd! dn PJ=0.00041 m=1 $X=3621760 $Y=80300 $D=8
D200 A5 vdd! dn PJ=0.0002 m=1 $X=3624020 $Y=13228100 $D=8
D201 A5 vdd! dn PJ=0.0002 m=1 $X=3624020 $Y=13438100 $D=8
D202 GND_PAD! VDD_PAD! dn PJ=0.00041 m=1 $X=3624260 $Y=80300 $D=8
D203 gnd! A5 dn PJ=0.0002 m=1 $X=3626340 $Y=13232500 $D=8
D204 gnd! A5 dn PJ=0.0002 m=1 $X=3626340 $Y=13442500 $D=8
D205 A5 vdd! dn PJ=0.0002 m=1 $X=3628660 $Y=13228100 $D=8
D206 A5 vdd! dn PJ=0.0002 m=1 $X=3628660 $Y=13438100 $D=8
D207 vdd! VDD_PAD! dn PJ=0.00041 m=1 $X=3629260 $Y=80300 $D=8
D208 gnd! A5 dn PJ=0.0001 m=1 $X=3630980 $Y=13332500 $D=8
D209 gnd! A5 dn PJ=0.0001 m=1 $X=3630980 $Y=13542500 $D=8
D210 VDD_PAD! vdd! dn PJ=0.00041 m=1 $X=3631760 $Y=80300 $D=8
D211 A5 vdd! dn PJ=0.0001 m=1 $X=3634160 $Y=13228100 $D=8
D212 A5 vdd! dn PJ=0.0001 m=1 $X=3634160 $Y=13438100 $D=8
D213 GND_PAD! VDD_PAD! dn PJ=0.00041 m=1 $X=3634260 $Y=80300 $D=8
D214 gnd! A5 dn PJ=0.0002 m=1 $X=3636480 $Y=13232500 $D=8
D215 gnd! A5 dn PJ=0.0002 m=1 $X=3636480 $Y=13442500 $D=8
D216 A5 vdd! dn PJ=0.0002 m=1 $X=3638800 $Y=13228100 $D=8
D217 A5 vdd! dn PJ=0.0002 m=1 $X=3638800 $Y=13438100 $D=8
D218 vdd! VDD_PAD! dn PJ=0.00041 m=1 $X=3639260 $Y=80300 $D=8
D219 gnd! A5 dn PJ=0.0002 m=1 $X=3641120 $Y=13232500 $D=8
D220 gnd! A5 dn PJ=0.0002 m=1 $X=3641120 $Y=13442500 $D=8
D221 VDD_PAD! vdd! dn PJ=0.00041 m=1 $X=3641760 $Y=80300 $D=8
D222 A5 vdd! dn PJ=0.0002 m=1 $X=3643440 $Y=13228100 $D=8
D223 A5 vdd! dn PJ=0.0002 m=1 $X=3643440 $Y=13438100 $D=8
D224 GND_PAD! VDD_PAD! dn PJ=0.00041 m=1 $X=3644260 $Y=80300 $D=8
D225 gnd! A5 dn PJ=0.0001 m=1 $X=3645760 $Y=13332500 $D=8
D226 gnd! A5 dn PJ=0.0001 m=1 $X=3645760 $Y=13542500 $D=8
D227 A5 vdd! dn PJ=0.0001 m=1 $X=3648940 $Y=13228100 $D=8
D228 A5 vdd! dn PJ=0.0001 m=1 $X=3648940 $Y=13438100 $D=8
D229 gnd! A5 dn PJ=0.0002 m=1 $X=3651260 $Y=13232500 $D=8
D230 gnd! A5 dn PJ=0.0002 m=1 $X=3651260 $Y=13442500 $D=8
D231 A5 vdd! dn PJ=0.0002 m=1 $X=3653580 $Y=13228100 $D=8
D232 A5 vdd! dn PJ=0.0002 m=1 $X=3653580 $Y=13438100 $D=8
D233 gnd! A5 dn PJ=0.0002 m=1 $X=3655900 $Y=13232500 $D=8
D234 gnd! A5 dn PJ=0.0002 m=1 $X=3655900 $Y=13442500 $D=8
D235 A5 vdd! dn PJ=0.0002 m=1 $X=3658220 $Y=13228100 $D=8
D236 A5 vdd! dn PJ=0.0002 m=1 $X=3658220 $Y=13438100 $D=8
D237 gnd! A5 dn PJ=0.0001 m=1 $X=3660540 $Y=13332500 $D=8
D238 gnd! A5 dn PJ=0.0001 m=1 $X=3660540 $Y=13542500 $D=8
D239 A5 vdd! dn PJ=0.0001 m=1 $X=3663720 $Y=13228100 $D=8
D240 A5 vdd! dn PJ=0.0001 m=1 $X=3663720 $Y=13438100 $D=8
D241 gnd! A5 dn PJ=0.0002 m=1 $X=3666040 $Y=13232500 $D=8
D242 gnd! A5 dn PJ=0.0002 m=1 $X=3666040 $Y=13442500 $D=8
D243 A5 vdd! dn PJ=0.0002 m=1 $X=3668360 $Y=13228100 $D=8
D244 A5 vdd! dn PJ=0.0002 m=1 $X=3668360 $Y=13438100 $D=8
D245 gnd! A5 dn PJ=0.0002 m=1 $X=3670680 $Y=13232500 $D=8
D246 gnd! A5 dn PJ=0.0002 m=1 $X=3670680 $Y=13442500 $D=8
D247 A5 vdd! dn PJ=0.0002 m=1 $X=3673000 $Y=13228100 $D=8
D248 A5 vdd! dn PJ=0.0002 m=1 $X=3673000 $Y=13438100 $D=8
D249 gnd! A5 dn PJ=0.0001 m=1 $X=3675320 $Y=13332500 $D=8
D250 gnd! A5 dn PJ=0.0001 m=1 $X=3675320 $Y=13542500 $D=8
D251 A5 vdd! dn PJ=0.0001 m=1 $X=3678500 $Y=13228100 $D=8
D252 A5 vdd! dn PJ=0.0001 m=1 $X=3678500 $Y=13438100 $D=8
D253 gnd! A5 dn PJ=0.0002 m=1 $X=3680820 $Y=13232500 $D=8
D254 gnd! A5 dn PJ=0.0002 m=1 $X=3680820 $Y=13442500 $D=8
D255 A5 vdd! dn PJ=0.0002 m=1 $X=3683140 $Y=13228100 $D=8
D256 A5 vdd! dn PJ=0.0002 m=1 $X=3683140 $Y=13438100 $D=8
D257 gnd! A5 dn PJ=0.0002 m=1 $X=3685460 $Y=13232500 $D=8
D258 gnd! A5 dn PJ=0.0002 m=1 $X=3685460 $Y=13442500 $D=8
D259 A5 vdd! dn PJ=0.0002 m=1 $X=3687780 $Y=13228100 $D=8
D260 A5 vdd! dn PJ=0.0002 m=1 $X=3687780 $Y=13438100 $D=8
D261 gnd! A5 dn PJ=0.0001 m=1 $X=3690100 $Y=13332500 $D=8
D262 gnd! A5 dn PJ=0.0001 m=1 $X=3690100 $Y=13542500 $D=8
D263 A5 vdd! dn PJ=0.0001 m=1 $X=3693280 $Y=13228100 $D=8
D264 A5 vdd! dn PJ=0.0001 m=1 $X=3693280 $Y=13438100 $D=8
D265 gnd! A5 dn PJ=0.0002 m=1 $X=3695600 $Y=13232500 $D=8
D266 gnd! A5 dn PJ=0.0002 m=1 $X=3695600 $Y=13442500 $D=8
D267 A5 vdd! dn PJ=0.0002 m=1 $X=3697920 $Y=13228100 $D=8
D268 A5 vdd! dn PJ=0.0002 m=1 $X=3697920 $Y=13438100 $D=8
D269 gnd! A5 dn PJ=0.0002 m=1 $X=3700240 $Y=13232500 $D=8
D270 gnd! A5 dn PJ=0.0002 m=1 $X=3700240 $Y=13442500 $D=8
D271 A5 vdd! dn PJ=0.0002 m=1 $X=3702560 $Y=13228100 $D=8
D272 A5 vdd! dn PJ=0.0002 m=1 $X=3702560 $Y=13438100 $D=8
D273 gnd! A5 dn PJ=0.0001 m=1 $X=3704880 $Y=13332500 $D=8
D274 gnd! A5 dn PJ=0.0001 m=1 $X=3704880 $Y=13542500 $D=8
D275 A5 vdd! dn PJ=0.0001 m=1 $X=3708060 $Y=13228100 $D=8
D276 A5 vdd! dn PJ=0.0001 m=1 $X=3708060 $Y=13438100 $D=8
D277 gnd! A5 dn PJ=0.0002 m=1 $X=3710380 $Y=13232500 $D=8
D278 gnd! A5 dn PJ=0.0002 m=1 $X=3710380 $Y=13442500 $D=8
D279 A5 vdd! dn PJ=0.0002 m=1 $X=3712700 $Y=13228100 $D=8
D280 A5 vdd! dn PJ=0.0002 m=1 $X=3712700 $Y=13438100 $D=8
D281 gnd! A5 dn PJ=0.0002 m=1 $X=3715020 $Y=13232500 $D=8
D282 gnd! A5 dn PJ=0.0002 m=1 $X=3715020 $Y=13442500 $D=8
D283 A8 vdd! dn PJ=0.0002 m=1 $X=5444020 $Y=13228100 $D=8
D284 A8 vdd! dn PJ=0.0002 m=1 $X=5444020 $Y=13438100 $D=8
D285 gnd! A8 dn PJ=0.0002 m=1 $X=5446340 $Y=13232500 $D=8
D286 gnd! A8 dn PJ=0.0002 m=1 $X=5446340 $Y=13442500 $D=8
D287 A8 vdd! dn PJ=0.0002 m=1 $X=5448660 $Y=13228100 $D=8
D288 A8 vdd! dn PJ=0.0002 m=1 $X=5448660 $Y=13438100 $D=8
D289 gnd! A8 dn PJ=0.0001 m=1 $X=5450980 $Y=13332500 $D=8
D290 gnd! A8 dn PJ=0.0001 m=1 $X=5450980 $Y=13542500 $D=8
D291 A8 vdd! dn PJ=0.0001 m=1 $X=5454160 $Y=13228100 $D=8
D292 A8 vdd! dn PJ=0.0001 m=1 $X=5454160 $Y=13438100 $D=8
D293 gnd! A8 dn PJ=0.0002 m=1 $X=5456480 $Y=13232500 $D=8
D294 gnd! A8 dn PJ=0.0002 m=1 $X=5456480 $Y=13442500 $D=8
D295 A8 vdd! dn PJ=0.0002 m=1 $X=5458800 $Y=13228100 $D=8
D296 A8 vdd! dn PJ=0.0002 m=1 $X=5458800 $Y=13438100 $D=8
D297 gnd! A8 dn PJ=0.0002 m=1 $X=5461120 $Y=13232500 $D=8
D298 gnd! A8 dn PJ=0.0002 m=1 $X=5461120 $Y=13442500 $D=8
D299 A8 vdd! dn PJ=0.0002 m=1 $X=5463440 $Y=13228100 $D=8
D300 A8 vdd! dn PJ=0.0002 m=1 $X=5463440 $Y=13438100 $D=8
D301 gnd! A8 dn PJ=0.0001 m=1 $X=5465760 $Y=13332500 $D=8
D302 gnd! A8 dn PJ=0.0001 m=1 $X=5465760 $Y=13542500 $D=8
D303 A8 vdd! dn PJ=0.0001 m=1 $X=5468940 $Y=13228100 $D=8
D304 A8 vdd! dn PJ=0.0001 m=1 $X=5468940 $Y=13438100 $D=8
D305 gnd! A8 dn PJ=0.0002 m=1 $X=5471260 $Y=13232500 $D=8
D306 gnd! A8 dn PJ=0.0002 m=1 $X=5471260 $Y=13442500 $D=8
D307 A8 vdd! dn PJ=0.0002 m=1 $X=5473580 $Y=13228100 $D=8
D308 A8 vdd! dn PJ=0.0002 m=1 $X=5473580 $Y=13438100 $D=8
D309 gnd! A8 dn PJ=0.0002 m=1 $X=5475900 $Y=13232500 $D=8
D310 gnd! A8 dn PJ=0.0002 m=1 $X=5475900 $Y=13442500 $D=8
D311 A8 vdd! dn PJ=0.0002 m=1 $X=5478220 $Y=13228100 $D=8
D312 A8 vdd! dn PJ=0.0002 m=1 $X=5478220 $Y=13438100 $D=8
D313 gnd! A8 dn PJ=0.0001 m=1 $X=5480540 $Y=13332500 $D=8
D314 gnd! A8 dn PJ=0.0001 m=1 $X=5480540 $Y=13542500 $D=8
D315 A8 vdd! dn PJ=0.0001 m=1 $X=5483720 $Y=13228100 $D=8
D316 A8 vdd! dn PJ=0.0001 m=1 $X=5483720 $Y=13438100 $D=8
D317 gnd! A8 dn PJ=0.0002 m=1 $X=5486040 $Y=13232500 $D=8
D318 gnd! A8 dn PJ=0.0002 m=1 $X=5486040 $Y=13442500 $D=8
D319 A8 vdd! dn PJ=0.0002 m=1 $X=5488360 $Y=13228100 $D=8
D320 A8 vdd! dn PJ=0.0002 m=1 $X=5488360 $Y=13438100 $D=8
D321 gnd! A8 dn PJ=0.0002 m=1 $X=5490680 $Y=13232500 $D=8
D322 gnd! A8 dn PJ=0.0002 m=1 $X=5490680 $Y=13442500 $D=8
D323 A8 vdd! dn PJ=0.0002 m=1 $X=5493000 $Y=13228100 $D=8
D324 A8 vdd! dn PJ=0.0002 m=1 $X=5493000 $Y=13438100 $D=8
D325 gnd! A8 dn PJ=0.0001 m=1 $X=5495320 $Y=13332500 $D=8
D326 gnd! A8 dn PJ=0.0001 m=1 $X=5495320 $Y=13542500 $D=8
D327 A8 vdd! dn PJ=0.0001 m=1 $X=5498500 $Y=13228100 $D=8
D328 A8 vdd! dn PJ=0.0001 m=1 $X=5498500 $Y=13438100 $D=8
D329 gnd! A8 dn PJ=0.0002 m=1 $X=5500820 $Y=13232500 $D=8
D330 gnd! A8 dn PJ=0.0002 m=1 $X=5500820 $Y=13442500 $D=8
D331 A8 vdd! dn PJ=0.0002 m=1 $X=5503140 $Y=13228100 $D=8
D332 A8 vdd! dn PJ=0.0002 m=1 $X=5503140 $Y=13438100 $D=8
D333 gnd! A8 dn PJ=0.0002 m=1 $X=5505460 $Y=13232500 $D=8
D334 gnd! A8 dn PJ=0.0002 m=1 $X=5505460 $Y=13442500 $D=8
D335 A8 vdd! dn PJ=0.0002 m=1 $X=5507780 $Y=13228100 $D=8
D336 A8 vdd! dn PJ=0.0002 m=1 $X=5507780 $Y=13438100 $D=8
D337 gnd! A8 dn PJ=0.0001 m=1 $X=5510100 $Y=13332500 $D=8
D338 gnd! A8 dn PJ=0.0001 m=1 $X=5510100 $Y=13542500 $D=8
D339 A8 vdd! dn PJ=0.0001 m=1 $X=5513280 $Y=13228100 $D=8
D340 A8 vdd! dn PJ=0.0001 m=1 $X=5513280 $Y=13438100 $D=8
D341 gnd! A8 dn PJ=0.0002 m=1 $X=5515600 $Y=13232500 $D=8
D342 gnd! A8 dn PJ=0.0002 m=1 $X=5515600 $Y=13442500 $D=8
D343 A8 vdd! dn PJ=0.0002 m=1 $X=5517920 $Y=13228100 $D=8
D344 A8 vdd! dn PJ=0.0002 m=1 $X=5517920 $Y=13438100 $D=8
D345 gnd! A8 dn PJ=0.0002 m=1 $X=5520240 $Y=13232500 $D=8
D346 gnd! A8 dn PJ=0.0002 m=1 $X=5520240 $Y=13442500 $D=8
D347 A8 vdd! dn PJ=0.0002 m=1 $X=5522560 $Y=13228100 $D=8
D348 A8 vdd! dn PJ=0.0002 m=1 $X=5522560 $Y=13438100 $D=8
D349 gnd! A8 dn PJ=0.0001 m=1 $X=5524880 $Y=13332500 $D=8
D350 gnd! A8 dn PJ=0.0001 m=1 $X=5524880 $Y=13542500 $D=8
D351 A8 vdd! dn PJ=0.0001 m=1 $X=5528060 $Y=13228100 $D=8
D352 A8 vdd! dn PJ=0.0001 m=1 $X=5528060 $Y=13438100 $D=8
D353 gnd! A8 dn PJ=0.0002 m=1 $X=5530380 $Y=13232500 $D=8
D354 gnd! A8 dn PJ=0.0002 m=1 $X=5530380 $Y=13442500 $D=8
D355 A8 vdd! dn PJ=0.0002 m=1 $X=5532700 $Y=13228100 $D=8
D356 A8 vdd! dn PJ=0.0002 m=1 $X=5532700 $Y=13438100 $D=8
D357 gnd! A8 dn PJ=0.0002 m=1 $X=5535020 $Y=13232500 $D=8
D358 gnd! A8 dn PJ=0.0002 m=1 $X=5535020 $Y=13442500 $D=8
D359 A9 vdd! dn PJ=0.0002 m=1 $X=5704020 $Y=13228100 $D=8
D360 A9 vdd! dn PJ=0.0002 m=1 $X=5704020 $Y=13438100 $D=8
D361 gnd! A9 dn PJ=0.0002 m=1 $X=5706340 $Y=13232500 $D=8
D362 gnd! A9 dn PJ=0.0002 m=1 $X=5706340 $Y=13442500 $D=8
D363 A9 vdd! dn PJ=0.0002 m=1 $X=5708660 $Y=13228100 $D=8
D364 A9 vdd! dn PJ=0.0002 m=1 $X=5708660 $Y=13438100 $D=8
D365 gnd! A9 dn PJ=0.0001 m=1 $X=5710980 $Y=13332500 $D=8
D366 gnd! A9 dn PJ=0.0001 m=1 $X=5710980 $Y=13542500 $D=8
D367 A9 vdd! dn PJ=0.0001 m=1 $X=5714160 $Y=13228100 $D=8
D368 A9 vdd! dn PJ=0.0001 m=1 $X=5714160 $Y=13438100 $D=8
D369 gnd! A9 dn PJ=0.0002 m=1 $X=5716480 $Y=13232500 $D=8
D370 gnd! A9 dn PJ=0.0002 m=1 $X=5716480 $Y=13442500 $D=8
D371 A9 vdd! dn PJ=0.0002 m=1 $X=5718800 $Y=13228100 $D=8
D372 A9 vdd! dn PJ=0.0002 m=1 $X=5718800 $Y=13438100 $D=8
D373 gnd! A9 dn PJ=0.0002 m=1 $X=5721120 $Y=13232500 $D=8
D374 gnd! A9 dn PJ=0.0002 m=1 $X=5721120 $Y=13442500 $D=8
D375 A9 vdd! dn PJ=0.0002 m=1 $X=5723440 $Y=13228100 $D=8
D376 A9 vdd! dn PJ=0.0002 m=1 $X=5723440 $Y=13438100 $D=8
D377 gnd! A9 dn PJ=0.0001 m=1 $X=5725760 $Y=13332500 $D=8
D378 gnd! A9 dn PJ=0.0001 m=1 $X=5725760 $Y=13542500 $D=8
D379 A9 vdd! dn PJ=0.0001 m=1 $X=5728940 $Y=13228100 $D=8
D380 A9 vdd! dn PJ=0.0001 m=1 $X=5728940 $Y=13438100 $D=8
D381 gnd! A9 dn PJ=0.0002 m=1 $X=5731260 $Y=13232500 $D=8
D382 gnd! A9 dn PJ=0.0002 m=1 $X=5731260 $Y=13442500 $D=8
D383 A9 vdd! dn PJ=0.0002 m=1 $X=5733580 $Y=13228100 $D=8
D384 A9 vdd! dn PJ=0.0002 m=1 $X=5733580 $Y=13438100 $D=8
D385 gnd! A9 dn PJ=0.0002 m=1 $X=5735900 $Y=13232500 $D=8
D386 gnd! A9 dn PJ=0.0002 m=1 $X=5735900 $Y=13442500 $D=8
D387 A9 vdd! dn PJ=0.0002 m=1 $X=5738220 $Y=13228100 $D=8
D388 A9 vdd! dn PJ=0.0002 m=1 $X=5738220 $Y=13438100 $D=8
D389 gnd! A9 dn PJ=0.0001 m=1 $X=5740540 $Y=13332500 $D=8
D390 gnd! A9 dn PJ=0.0001 m=1 $X=5740540 $Y=13542500 $D=8
D391 A9 vdd! dn PJ=0.0001 m=1 $X=5743720 $Y=13228100 $D=8
D392 A9 vdd! dn PJ=0.0001 m=1 $X=5743720 $Y=13438100 $D=8
D393 gnd! A9 dn PJ=0.0002 m=1 $X=5746040 $Y=13232500 $D=8
D394 gnd! A9 dn PJ=0.0002 m=1 $X=5746040 $Y=13442500 $D=8
D395 A9 vdd! dn PJ=0.0002 m=1 $X=5748360 $Y=13228100 $D=8
D396 A9 vdd! dn PJ=0.0002 m=1 $X=5748360 $Y=13438100 $D=8
D397 gnd! A9 dn PJ=0.0002 m=1 $X=5750680 $Y=13232500 $D=8
D398 gnd! A9 dn PJ=0.0002 m=1 $X=5750680 $Y=13442500 $D=8
D399 A9 vdd! dn PJ=0.0002 m=1 $X=5753000 $Y=13228100 $D=8
D400 A9 vdd! dn PJ=0.0002 m=1 $X=5753000 $Y=13438100 $D=8
D401 gnd! A9 dn PJ=0.0001 m=1 $X=5755320 $Y=13332500 $D=8
D402 gnd! A9 dn PJ=0.0001 m=1 $X=5755320 $Y=13542500 $D=8
D403 A9 vdd! dn PJ=0.0001 m=1 $X=5758500 $Y=13228100 $D=8
D404 A9 vdd! dn PJ=0.0001 m=1 $X=5758500 $Y=13438100 $D=8
D405 gnd! A9 dn PJ=0.0002 m=1 $X=5760820 $Y=13232500 $D=8
D406 gnd! A9 dn PJ=0.0002 m=1 $X=5760820 $Y=13442500 $D=8
D407 A9 vdd! dn PJ=0.0002 m=1 $X=5763140 $Y=13228100 $D=8
D408 A9 vdd! dn PJ=0.0002 m=1 $X=5763140 $Y=13438100 $D=8
D409 gnd! A9 dn PJ=0.0002 m=1 $X=5765460 $Y=13232500 $D=8
D410 gnd! A9 dn PJ=0.0002 m=1 $X=5765460 $Y=13442500 $D=8
D411 A9 vdd! dn PJ=0.0002 m=1 $X=5767780 $Y=13228100 $D=8
D412 A9 vdd! dn PJ=0.0002 m=1 $X=5767780 $Y=13438100 $D=8
D413 gnd! A9 dn PJ=0.0001 m=1 $X=5770100 $Y=13332500 $D=8
D414 gnd! A9 dn PJ=0.0001 m=1 $X=5770100 $Y=13542500 $D=8
D415 A9 vdd! dn PJ=0.0001 m=1 $X=5773280 $Y=13228100 $D=8
D416 A9 vdd! dn PJ=0.0001 m=1 $X=5773280 $Y=13438100 $D=8
D417 gnd! A9 dn PJ=0.0002 m=1 $X=5775600 $Y=13232500 $D=8
D418 gnd! A9 dn PJ=0.0002 m=1 $X=5775600 $Y=13442500 $D=8
D419 A9 vdd! dn PJ=0.0002 m=1 $X=5777920 $Y=13228100 $D=8
D420 A9 vdd! dn PJ=0.0002 m=1 $X=5777920 $Y=13438100 $D=8
D421 gnd! A9 dn PJ=0.0002 m=1 $X=5780240 $Y=13232500 $D=8
D422 gnd! A9 dn PJ=0.0002 m=1 $X=5780240 $Y=13442500 $D=8
D423 A9 vdd! dn PJ=0.0002 m=1 $X=5782560 $Y=13228100 $D=8
D424 A9 vdd! dn PJ=0.0002 m=1 $X=5782560 $Y=13438100 $D=8
D425 gnd! A9 dn PJ=0.0001 m=1 $X=5784880 $Y=13332500 $D=8
D426 gnd! A9 dn PJ=0.0001 m=1 $X=5784880 $Y=13542500 $D=8
D427 A9 vdd! dn PJ=0.0001 m=1 $X=5788060 $Y=13228100 $D=8
D428 A9 vdd! dn PJ=0.0001 m=1 $X=5788060 $Y=13438100 $D=8
D429 gnd! A9 dn PJ=0.0002 m=1 $X=5790380 $Y=13232500 $D=8
D430 gnd! A9 dn PJ=0.0002 m=1 $X=5790380 $Y=13442500 $D=8
D431 A9 vdd! dn PJ=0.0002 m=1 $X=5792700 $Y=13228100 $D=8
D432 A9 vdd! dn PJ=0.0002 m=1 $X=5792700 $Y=13438100 $D=8
D433 gnd! A9 dn PJ=0.0002 m=1 $X=5795020 $Y=13232500 $D=8
D434 gnd! A9 dn PJ=0.0002 m=1 $X=5795020 $Y=13442500 $D=8
D435 A10 vdd! dn PJ=0.0002 m=1 $X=5964020 $Y=13228100 $D=8
D436 A10 vdd! dn PJ=0.0002 m=1 $X=5964020 $Y=13438100 $D=8
D437 gnd! A10 dn PJ=0.0002 m=1 $X=5966340 $Y=13232500 $D=8
D438 gnd! A10 dn PJ=0.0002 m=1 $X=5966340 $Y=13442500 $D=8
D439 A10 vdd! dn PJ=0.0002 m=1 $X=5968660 $Y=13228100 $D=8
D440 A10 vdd! dn PJ=0.0002 m=1 $X=5968660 $Y=13438100 $D=8
D441 gnd! A10 dn PJ=0.0001 m=1 $X=5970980 $Y=13332500 $D=8
D442 gnd! A10 dn PJ=0.0001 m=1 $X=5970980 $Y=13542500 $D=8
D443 A10 vdd! dn PJ=0.0001 m=1 $X=5974160 $Y=13228100 $D=8
D444 A10 vdd! dn PJ=0.0001 m=1 $X=5974160 $Y=13438100 $D=8
D445 gnd! A10 dn PJ=0.0002 m=1 $X=5976480 $Y=13232500 $D=8
D446 gnd! A10 dn PJ=0.0002 m=1 $X=5976480 $Y=13442500 $D=8
D447 A10 vdd! dn PJ=0.0002 m=1 $X=5978800 $Y=13228100 $D=8
D448 A10 vdd! dn PJ=0.0002 m=1 $X=5978800 $Y=13438100 $D=8
D449 gnd! A10 dn PJ=0.0002 m=1 $X=5981120 $Y=13232500 $D=8
D450 gnd! A10 dn PJ=0.0002 m=1 $X=5981120 $Y=13442500 $D=8
D451 A10 vdd! dn PJ=0.0002 m=1 $X=5983440 $Y=13228100 $D=8
D452 A10 vdd! dn PJ=0.0002 m=1 $X=5983440 $Y=13438100 $D=8
D453 gnd! A10 dn PJ=0.0001 m=1 $X=5985760 $Y=13332500 $D=8
D454 gnd! A10 dn PJ=0.0001 m=1 $X=5985760 $Y=13542500 $D=8
D455 A10 vdd! dn PJ=0.0001 m=1 $X=5988940 $Y=13228100 $D=8
D456 A10 vdd! dn PJ=0.0001 m=1 $X=5988940 $Y=13438100 $D=8
D457 gnd! A10 dn PJ=0.0002 m=1 $X=5991260 $Y=13232500 $D=8
D458 gnd! A10 dn PJ=0.0002 m=1 $X=5991260 $Y=13442500 $D=8
D459 A10 vdd! dn PJ=0.0002 m=1 $X=5993580 $Y=13228100 $D=8
D460 A10 vdd! dn PJ=0.0002 m=1 $X=5993580 $Y=13438100 $D=8
D461 gnd! A10 dn PJ=0.0002 m=1 $X=5995900 $Y=13232500 $D=8
D462 gnd! A10 dn PJ=0.0002 m=1 $X=5995900 $Y=13442500 $D=8
D463 A10 vdd! dn PJ=0.0002 m=1 $X=5998220 $Y=13228100 $D=8
D464 A10 vdd! dn PJ=0.0002 m=1 $X=5998220 $Y=13438100 $D=8
D465 gnd! A10 dn PJ=0.0001 m=1 $X=6000540 $Y=13332500 $D=8
D466 gnd! A10 dn PJ=0.0001 m=1 $X=6000540 $Y=13542500 $D=8
D467 A10 vdd! dn PJ=0.0001 m=1 $X=6003720 $Y=13228100 $D=8
D468 A10 vdd! dn PJ=0.0001 m=1 $X=6003720 $Y=13438100 $D=8
D469 gnd! A10 dn PJ=0.0002 m=1 $X=6006040 $Y=13232500 $D=8
D470 gnd! A10 dn PJ=0.0002 m=1 $X=6006040 $Y=13442500 $D=8
D471 A10 vdd! dn PJ=0.0002 m=1 $X=6008360 $Y=13228100 $D=8
D472 A10 vdd! dn PJ=0.0002 m=1 $X=6008360 $Y=13438100 $D=8
D473 gnd! A10 dn PJ=0.0002 m=1 $X=6010680 $Y=13232500 $D=8
D474 gnd! A10 dn PJ=0.0002 m=1 $X=6010680 $Y=13442500 $D=8
D475 A10 vdd! dn PJ=0.0002 m=1 $X=6013000 $Y=13228100 $D=8
D476 A10 vdd! dn PJ=0.0002 m=1 $X=6013000 $Y=13438100 $D=8
D477 gnd! A10 dn PJ=0.0001 m=1 $X=6015320 $Y=13332500 $D=8
D478 gnd! A10 dn PJ=0.0001 m=1 $X=6015320 $Y=13542500 $D=8
D479 A10 vdd! dn PJ=0.0001 m=1 $X=6018500 $Y=13228100 $D=8
D480 A10 vdd! dn PJ=0.0001 m=1 $X=6018500 $Y=13438100 $D=8
D481 gnd! A10 dn PJ=0.0002 m=1 $X=6020820 $Y=13232500 $D=8
D482 gnd! A10 dn PJ=0.0002 m=1 $X=6020820 $Y=13442500 $D=8
D483 A10 vdd! dn PJ=0.0002 m=1 $X=6023140 $Y=13228100 $D=8
D484 A10 vdd! dn PJ=0.0002 m=1 $X=6023140 $Y=13438100 $D=8
D485 gnd! A10 dn PJ=0.0002 m=1 $X=6025460 $Y=13232500 $D=8
D486 gnd! A10 dn PJ=0.0002 m=1 $X=6025460 $Y=13442500 $D=8
D487 A10 vdd! dn PJ=0.0002 m=1 $X=6027780 $Y=13228100 $D=8
D488 A10 vdd! dn PJ=0.0002 m=1 $X=6027780 $Y=13438100 $D=8
D489 gnd! A10 dn PJ=0.0001 m=1 $X=6030100 $Y=13332500 $D=8
D490 gnd! A10 dn PJ=0.0001 m=1 $X=6030100 $Y=13542500 $D=8
D491 A10 vdd! dn PJ=0.0001 m=1 $X=6033280 $Y=13228100 $D=8
D492 A10 vdd! dn PJ=0.0001 m=1 $X=6033280 $Y=13438100 $D=8
D493 gnd! A10 dn PJ=0.0002 m=1 $X=6035600 $Y=13232500 $D=8
D494 gnd! A10 dn PJ=0.0002 m=1 $X=6035600 $Y=13442500 $D=8
D495 A10 vdd! dn PJ=0.0002 m=1 $X=6037920 $Y=13228100 $D=8
D496 A10 vdd! dn PJ=0.0002 m=1 $X=6037920 $Y=13438100 $D=8
D497 gnd! A10 dn PJ=0.0002 m=1 $X=6040240 $Y=13232500 $D=8
D498 gnd! A10 dn PJ=0.0002 m=1 $X=6040240 $Y=13442500 $D=8
D499 A10 vdd! dn PJ=0.0002 m=1 $X=6042560 $Y=13228100 $D=8
D500 A10 vdd! dn PJ=0.0002 m=1 $X=6042560 $Y=13438100 $D=8
D501 gnd! A10 dn PJ=0.0001 m=1 $X=6044880 $Y=13332500 $D=8
D502 gnd! A10 dn PJ=0.0001 m=1 $X=6044880 $Y=13542500 $D=8
D503 A10 vdd! dn PJ=0.0001 m=1 $X=6048060 $Y=13228100 $D=8
D504 A10 vdd! dn PJ=0.0001 m=1 $X=6048060 $Y=13438100 $D=8
D505 gnd! A10 dn PJ=0.0002 m=1 $X=6050380 $Y=13232500 $D=8
D506 gnd! A10 dn PJ=0.0002 m=1 $X=6050380 $Y=13442500 $D=8
D507 A10 vdd! dn PJ=0.0002 m=1 $X=6052700 $Y=13228100 $D=8
D508 A10 vdd! dn PJ=0.0002 m=1 $X=6052700 $Y=13438100 $D=8
D509 gnd! A10 dn PJ=0.0002 m=1 $X=6055020 $Y=13232500 $D=8
D510 gnd! A10 dn PJ=0.0002 m=1 $X=6055020 $Y=13442500 $D=8
D511 CS1 vdd! dn PJ=0.0002 m=1 $X=6484020 $Y=13228100 $D=8
D512 CS1 vdd! dn PJ=0.0002 m=1 $X=6484020 $Y=13438100 $D=8
D513 gnd! CS1 dn PJ=0.0002 m=1 $X=6486340 $Y=13232500 $D=8
D514 gnd! CS1 dn PJ=0.0002 m=1 $X=6486340 $Y=13442500 $D=8
D515 CS1 vdd! dn PJ=0.0002 m=1 $X=6488660 $Y=13228100 $D=8
D516 CS1 vdd! dn PJ=0.0002 m=1 $X=6488660 $Y=13438100 $D=8
D517 gnd! CS1 dn PJ=0.0001 m=1 $X=6490980 $Y=13332500 $D=8
D518 gnd! CS1 dn PJ=0.0001 m=1 $X=6490980 $Y=13542500 $D=8
D519 CS1 vdd! dn PJ=0.0001 m=1 $X=6494160 $Y=13228100 $D=8
D520 CS1 vdd! dn PJ=0.0001 m=1 $X=6494160 $Y=13438100 $D=8
D521 gnd! CS1 dn PJ=0.0002 m=1 $X=6496480 $Y=13232500 $D=8
D522 gnd! CS1 dn PJ=0.0002 m=1 $X=6496480 $Y=13442500 $D=8
D523 CS1 vdd! dn PJ=0.0002 m=1 $X=6498800 $Y=13228100 $D=8
D524 CS1 vdd! dn PJ=0.0002 m=1 $X=6498800 $Y=13438100 $D=8
D525 gnd! CS1 dn PJ=0.0002 m=1 $X=6501120 $Y=13232500 $D=8
D526 gnd! CS1 dn PJ=0.0002 m=1 $X=6501120 $Y=13442500 $D=8
D527 CS1 vdd! dn PJ=0.0002 m=1 $X=6503440 $Y=13228100 $D=8
D528 CS1 vdd! dn PJ=0.0002 m=1 $X=6503440 $Y=13438100 $D=8
D529 gnd! CS1 dn PJ=0.0001 m=1 $X=6505760 $Y=13332500 $D=8
D530 gnd! CS1 dn PJ=0.0001 m=1 $X=6505760 $Y=13542500 $D=8
D531 CS1 vdd! dn PJ=0.0001 m=1 $X=6508940 $Y=13228100 $D=8
D532 CS1 vdd! dn PJ=0.0001 m=1 $X=6508940 $Y=13438100 $D=8
D533 gnd! CS1 dn PJ=0.0002 m=1 $X=6511260 $Y=13232500 $D=8
D534 gnd! CS1 dn PJ=0.0002 m=1 $X=6511260 $Y=13442500 $D=8
D535 CS1 vdd! dn PJ=0.0002 m=1 $X=6513580 $Y=13228100 $D=8
D536 CS1 vdd! dn PJ=0.0002 m=1 $X=6513580 $Y=13438100 $D=8
D537 gnd! CS1 dn PJ=0.0002 m=1 $X=6515900 $Y=13232500 $D=8
D538 gnd! CS1 dn PJ=0.0002 m=1 $X=6515900 $Y=13442500 $D=8
D539 CS1 vdd! dn PJ=0.0002 m=1 $X=6518220 $Y=13228100 $D=8
D540 CS1 vdd! dn PJ=0.0002 m=1 $X=6518220 $Y=13438100 $D=8
D541 gnd! CS1 dn PJ=0.0001 m=1 $X=6520540 $Y=13332500 $D=8
D542 gnd! CS1 dn PJ=0.0001 m=1 $X=6520540 $Y=13542500 $D=8
D543 CS1 vdd! dn PJ=0.0001 m=1 $X=6523720 $Y=13228100 $D=8
D544 CS1 vdd! dn PJ=0.0001 m=1 $X=6523720 $Y=13438100 $D=8
D545 gnd! CS1 dn PJ=0.0002 m=1 $X=6526040 $Y=13232500 $D=8
D546 gnd! CS1 dn PJ=0.0002 m=1 $X=6526040 $Y=13442500 $D=8
D547 CS1 vdd! dn PJ=0.0002 m=1 $X=6528360 $Y=13228100 $D=8
D548 CS1 vdd! dn PJ=0.0002 m=1 $X=6528360 $Y=13438100 $D=8
D549 gnd! CS1 dn PJ=0.0002 m=1 $X=6530680 $Y=13232500 $D=8
D550 gnd! CS1 dn PJ=0.0002 m=1 $X=6530680 $Y=13442500 $D=8
D551 CS1 vdd! dn PJ=0.0002 m=1 $X=6533000 $Y=13228100 $D=8
D552 CS1 vdd! dn PJ=0.0002 m=1 $X=6533000 $Y=13438100 $D=8
D553 gnd! CS1 dn PJ=0.0001 m=1 $X=6535320 $Y=13332500 $D=8
D554 gnd! CS1 dn PJ=0.0001 m=1 $X=6535320 $Y=13542500 $D=8
D555 CS1 vdd! dn PJ=0.0001 m=1 $X=6538500 $Y=13228100 $D=8
D556 CS1 vdd! dn PJ=0.0001 m=1 $X=6538500 $Y=13438100 $D=8
D557 gnd! CS1 dn PJ=0.0002 m=1 $X=6540820 $Y=13232500 $D=8
D558 gnd! CS1 dn PJ=0.0002 m=1 $X=6540820 $Y=13442500 $D=8
D559 CS1 vdd! dn PJ=0.0002 m=1 $X=6543140 $Y=13228100 $D=8
D560 CS1 vdd! dn PJ=0.0002 m=1 $X=6543140 $Y=13438100 $D=8
D561 gnd! CS1 dn PJ=0.0002 m=1 $X=6545460 $Y=13232500 $D=8
D562 gnd! CS1 dn PJ=0.0002 m=1 $X=6545460 $Y=13442500 $D=8
D563 CS1 vdd! dn PJ=0.0002 m=1 $X=6547780 $Y=13228100 $D=8
D564 CS1 vdd! dn PJ=0.0002 m=1 $X=6547780 $Y=13438100 $D=8
D565 gnd! CS1 dn PJ=0.0001 m=1 $X=6550100 $Y=13332500 $D=8
D566 gnd! CS1 dn PJ=0.0001 m=1 $X=6550100 $Y=13542500 $D=8
D567 CS1 vdd! dn PJ=0.0001 m=1 $X=6553280 $Y=13228100 $D=8
D568 CS1 vdd! dn PJ=0.0001 m=1 $X=6553280 $Y=13438100 $D=8
D569 gnd! CS1 dn PJ=0.0002 m=1 $X=6555600 $Y=13232500 $D=8
D570 gnd! CS1 dn PJ=0.0002 m=1 $X=6555600 $Y=13442500 $D=8
D571 CS1 vdd! dn PJ=0.0002 m=1 $X=6557920 $Y=13228100 $D=8
D572 CS1 vdd! dn PJ=0.0002 m=1 $X=6557920 $Y=13438100 $D=8
D573 gnd! CS1 dn PJ=0.0002 m=1 $X=6560240 $Y=13232500 $D=8
D574 gnd! CS1 dn PJ=0.0002 m=1 $X=6560240 $Y=13442500 $D=8
D575 CS1 vdd! dn PJ=0.0002 m=1 $X=6562560 $Y=13228100 $D=8
D576 CS1 vdd! dn PJ=0.0002 m=1 $X=6562560 $Y=13438100 $D=8
D577 gnd! CS1 dn PJ=0.0001 m=1 $X=6564880 $Y=13332500 $D=8
D578 gnd! CS1 dn PJ=0.0001 m=1 $X=6564880 $Y=13542500 $D=8
D579 CS1 vdd! dn PJ=0.0001 m=1 $X=6568060 $Y=13228100 $D=8
D580 CS1 vdd! dn PJ=0.0001 m=1 $X=6568060 $Y=13438100 $D=8
D581 gnd! CS1 dn PJ=0.0002 m=1 $X=6570380 $Y=13232500 $D=8
D582 gnd! CS1 dn PJ=0.0002 m=1 $X=6570380 $Y=13442500 $D=8
D583 CS1 vdd! dn PJ=0.0002 m=1 $X=6572700 $Y=13228100 $D=8
D584 CS1 vdd! dn PJ=0.0002 m=1 $X=6572700 $Y=13438100 $D=8
D585 gnd! CS1 dn PJ=0.0002 m=1 $X=6575020 $Y=13232500 $D=8
D586 gnd! CS1 dn PJ=0.0002 m=1 $X=6575020 $Y=13442500 $D=8
D587 vdd! VDD_PAD! dn PJ=0.00041 m=1 $X=7159060 $Y=80300 $D=8
D588 gnd! vdd! dn PJ=0.00041 m=1 $X=7161560 $Y=80300 $D=8
D589 vdd! VDD_PAD! dn PJ=0.00041 m=1 $X=7169060 $Y=80300 $D=8
D590 gnd! vdd! dn PJ=0.00041 m=1 $X=7171560 $Y=80300 $D=8
D591 vdd! VDD_PAD! dn PJ=0.00041 m=1 $X=7179060 $Y=80300 $D=8
D592 gnd! vdd! dn PJ=0.00041 m=1 $X=7181560 $Y=80300 $D=8
D593 vdd! VDD_PAD! dn PJ=0.00041 m=1 $X=7189060 $Y=80300 $D=8
D594 gnd! vdd! dn PJ=0.00041 m=1 $X=7191560 $Y=80300 $D=8
D595 vdd! VDD_PAD! dn PJ=0.00041 m=1 $X=7199060 $Y=80300 $D=8
D596 gnd! vdd! dn PJ=0.00041 m=1 $X=7201560 $Y=80300 $D=8
D597 vdd! VDD_PAD! dn PJ=0.00041 m=1 $X=7209060 $Y=80300 $D=8
D598 gnd! vdd! dn PJ=0.00041 m=1 $X=7211560 $Y=80300 $D=8
D599 vdd! VDD_PAD! dn PJ=0.00041 m=1 $X=7219060 $Y=80300 $D=8
D600 gnd! vdd! dn PJ=0.00041 m=1 $X=7221560 $Y=80300 $D=8
D601 vdd! VDD_PAD! dn PJ=0.00041 m=1 $X=7229060 $Y=80300 $D=8
D602 gnd! vdd! dn PJ=0.00041 m=1 $X=7231560 $Y=80300 $D=8
D603 vdd! VDD_PAD! dn PJ=0.00041 m=1 $X=7239060 $Y=80300 $D=8
D604 gnd! vdd! dn PJ=0.00041 m=1 $X=7241560 $Y=80300 $D=8
D605 gnd! vdd! dn PJ=0.00041 m=1 $X=7454280 $Y=80300 $D=8
D606 vdd! VDD_PAD! dn PJ=0.00041 m=1 $X=7461780 $Y=80300 $D=8
D607 gnd! vdd! dn PJ=0.00041 m=1 $X=7464280 $Y=80300 $D=8
D608 vdd! VDD_PAD! dn PJ=0.00041 m=1 $X=7471780 $Y=80300 $D=8
D609 gnd! vdd! dn PJ=0.00041 m=1 $X=7474280 $Y=80300 $D=8
D610 vdd! VDD_PAD! dn PJ=0.00041 m=1 $X=7481780 $Y=80300 $D=8
D611 gnd! vdd! dn PJ=0.00041 m=1 $X=7484280 $Y=80300 $D=8
D612 vdd! VDD_PAD! dn PJ=0.00041 m=1 $X=7491780 $Y=80300 $D=8
D613 gnd! vdd! dn PJ=0.00041 m=1 $X=7494280 $Y=80300 $D=8
D614 vdd! VDD_PAD! dn PJ=0.00041 m=1 $X=7501780 $Y=80300 $D=8
D615 gnd! vdd! dn PJ=0.00041 m=1 $X=7504280 $Y=80300 $D=8
D616 vdd! VDD_PAD! dn PJ=0.00041 m=1 $X=7511780 $Y=80300 $D=8
D617 gnd! vdd! dn PJ=0.00041 m=1 $X=7514280 $Y=80300 $D=8
D618 vdd! VDD_PAD! dn PJ=0.00041 m=1 $X=7521780 $Y=80300 $D=8
D619 A11 vdd! dn PJ=0.0002 m=1 $X=7524020 $Y=13228100 $D=8
D620 A11 vdd! dn PJ=0.0002 m=1 $X=7524020 $Y=13438100 $D=8
D621 gnd! vdd! dn PJ=0.00041 m=1 $X=7524280 $Y=80300 $D=8
D622 gnd! A11 dn PJ=0.0002 m=1 $X=7526340 $Y=13232500 $D=8
D623 gnd! A11 dn PJ=0.0002 m=1 $X=7526340 $Y=13442500 $D=8
D624 A11 vdd! dn PJ=0.0002 m=1 $X=7528660 $Y=13228100 $D=8
D625 A11 vdd! dn PJ=0.0002 m=1 $X=7528660 $Y=13438100 $D=8
D626 gnd! A11 dn PJ=0.0001 m=1 $X=7530980 $Y=13332500 $D=8
D627 gnd! A11 dn PJ=0.0001 m=1 $X=7530980 $Y=13542500 $D=8
D628 vdd! VDD_PAD! dn PJ=0.00041 m=1 $X=7531780 $Y=80300 $D=8
D629 A11 vdd! dn PJ=0.0001 m=1 $X=7534160 $Y=13228100 $D=8
D630 A11 vdd! dn PJ=0.0001 m=1 $X=7534160 $Y=13438100 $D=8
D631 gnd! vdd! dn PJ=0.00041 m=1 $X=7534280 $Y=80300 $D=8
D632 gnd! A11 dn PJ=0.0002 m=1 $X=7536480 $Y=13232500 $D=8
D633 gnd! A11 dn PJ=0.0002 m=1 $X=7536480 $Y=13442500 $D=8
D634 A11 vdd! dn PJ=0.0002 m=1 $X=7538800 $Y=13228100 $D=8
D635 A11 vdd! dn PJ=0.0002 m=1 $X=7538800 $Y=13438100 $D=8
D636 gnd! A11 dn PJ=0.0002 m=1 $X=7541120 $Y=13232500 $D=8
D637 gnd! A11 dn PJ=0.0002 m=1 $X=7541120 $Y=13442500 $D=8
D638 vdd! VDD_PAD! dn PJ=0.00041 m=1 $X=7541780 $Y=80300 $D=8
D639 A11 vdd! dn PJ=0.0002 m=1 $X=7543440 $Y=13228100 $D=8
D640 A11 vdd! dn PJ=0.0002 m=1 $X=7543440 $Y=13438100 $D=8
D641 gnd! vdd! dn PJ=0.00041 m=1 $X=7544280 $Y=80300 $D=8
D642 gnd! A11 dn PJ=0.0001 m=1 $X=7545760 $Y=13332500 $D=8
D643 gnd! A11 dn PJ=0.0001 m=1 $X=7545760 $Y=13542500 $D=8
D644 A11 vdd! dn PJ=0.0001 m=1 $X=7548940 $Y=13228100 $D=8
D645 A11 vdd! dn PJ=0.0001 m=1 $X=7548940 $Y=13438100 $D=8
D646 gnd! A11 dn PJ=0.0002 m=1 $X=7551260 $Y=13232500 $D=8
D647 gnd! A11 dn PJ=0.0002 m=1 $X=7551260 $Y=13442500 $D=8
D648 A11 vdd! dn PJ=0.0002 m=1 $X=7553580 $Y=13228100 $D=8
D649 A11 vdd! dn PJ=0.0002 m=1 $X=7553580 $Y=13438100 $D=8
D650 gnd! A11 dn PJ=0.0002 m=1 $X=7555900 $Y=13232500 $D=8
D651 gnd! A11 dn PJ=0.0002 m=1 $X=7555900 $Y=13442500 $D=8
D652 A11 vdd! dn PJ=0.0002 m=1 $X=7558220 $Y=13228100 $D=8
D653 A11 vdd! dn PJ=0.0002 m=1 $X=7558220 $Y=13438100 $D=8
D654 gnd! A11 dn PJ=0.0001 m=1 $X=7560540 $Y=13332500 $D=8
D655 gnd! A11 dn PJ=0.0001 m=1 $X=7560540 $Y=13542500 $D=8
D656 A11 vdd! dn PJ=0.0001 m=1 $X=7563720 $Y=13228100 $D=8
D657 A11 vdd! dn PJ=0.0001 m=1 $X=7563720 $Y=13438100 $D=8
D658 gnd! A11 dn PJ=0.0002 m=1 $X=7566040 $Y=13232500 $D=8
D659 gnd! A11 dn PJ=0.0002 m=1 $X=7566040 $Y=13442500 $D=8
D660 A11 vdd! dn PJ=0.0002 m=1 $X=7568360 $Y=13228100 $D=8
D661 A11 vdd! dn PJ=0.0002 m=1 $X=7568360 $Y=13438100 $D=8
D662 gnd! A11 dn PJ=0.0002 m=1 $X=7570680 $Y=13232500 $D=8
D663 gnd! A11 dn PJ=0.0002 m=1 $X=7570680 $Y=13442500 $D=8
D664 A11 vdd! dn PJ=0.0002 m=1 $X=7573000 $Y=13228100 $D=8
D665 A11 vdd! dn PJ=0.0002 m=1 $X=7573000 $Y=13438100 $D=8
D666 gnd! A11 dn PJ=0.0001 m=1 $X=7575320 $Y=13332500 $D=8
D667 gnd! A11 dn PJ=0.0001 m=1 $X=7575320 $Y=13542500 $D=8
D668 A11 vdd! dn PJ=0.0001 m=1 $X=7578500 $Y=13228100 $D=8
D669 A11 vdd! dn PJ=0.0001 m=1 $X=7578500 $Y=13438100 $D=8
D670 gnd! A11 dn PJ=0.0002 m=1 $X=7580820 $Y=13232500 $D=8
D671 gnd! A11 dn PJ=0.0002 m=1 $X=7580820 $Y=13442500 $D=8
D672 A11 vdd! dn PJ=0.0002 m=1 $X=7583140 $Y=13228100 $D=8
D673 A11 vdd! dn PJ=0.0002 m=1 $X=7583140 $Y=13438100 $D=8
D674 gnd! A11 dn PJ=0.0002 m=1 $X=7585460 $Y=13232500 $D=8
D675 gnd! A11 dn PJ=0.0002 m=1 $X=7585460 $Y=13442500 $D=8
D676 A11 vdd! dn PJ=0.0002 m=1 $X=7587780 $Y=13228100 $D=8
D677 A11 vdd! dn PJ=0.0002 m=1 $X=7587780 $Y=13438100 $D=8
D678 gnd! A11 dn PJ=0.0001 m=1 $X=7590100 $Y=13332500 $D=8
D679 gnd! A11 dn PJ=0.0001 m=1 $X=7590100 $Y=13542500 $D=8
D680 A11 vdd! dn PJ=0.0001 m=1 $X=7593280 $Y=13228100 $D=8
D681 A11 vdd! dn PJ=0.0001 m=1 $X=7593280 $Y=13438100 $D=8
D682 gnd! A11 dn PJ=0.0002 m=1 $X=7595600 $Y=13232500 $D=8
D683 gnd! A11 dn PJ=0.0002 m=1 $X=7595600 $Y=13442500 $D=8
D684 A11 vdd! dn PJ=0.0002 m=1 $X=7597920 $Y=13228100 $D=8
D685 A11 vdd! dn PJ=0.0002 m=1 $X=7597920 $Y=13438100 $D=8
D686 gnd! A11 dn PJ=0.0002 m=1 $X=7600240 $Y=13232500 $D=8
D687 gnd! A11 dn PJ=0.0002 m=1 $X=7600240 $Y=13442500 $D=8
D688 A11 vdd! dn PJ=0.0002 m=1 $X=7602560 $Y=13228100 $D=8
D689 A11 vdd! dn PJ=0.0002 m=1 $X=7602560 $Y=13438100 $D=8
D690 gnd! A11 dn PJ=0.0001 m=1 $X=7604880 $Y=13332500 $D=8
D691 gnd! A11 dn PJ=0.0001 m=1 $X=7604880 $Y=13542500 $D=8
D692 A11 vdd! dn PJ=0.0001 m=1 $X=7608060 $Y=13228100 $D=8
D693 A11 vdd! dn PJ=0.0001 m=1 $X=7608060 $Y=13438100 $D=8
D694 gnd! A11 dn PJ=0.0002 m=1 $X=7610380 $Y=13232500 $D=8
D695 gnd! A11 dn PJ=0.0002 m=1 $X=7610380 $Y=13442500 $D=8
D696 A11 vdd! dn PJ=0.0002 m=1 $X=7612700 $Y=13228100 $D=8
D697 A11 vdd! dn PJ=0.0002 m=1 $X=7612700 $Y=13438100 $D=8
D698 gnd! A11 dn PJ=0.0002 m=1 $X=7615020 $Y=13232500 $D=8
D699 gnd! A11 dn PJ=0.0002 m=1 $X=7615020 $Y=13442500 $D=8
D700 GND_PAD! VDD_PAD! dn PJ=0.00041 m=1 $X=7761540 $Y=80300 $D=8
D701 GND_PAD! VDD_PAD! dn PJ=0.00041 m=1 $X=7771540 $Y=80300 $D=8
D702 GND_PAD! VDD_PAD! dn PJ=0.00041 m=1 $X=7781540 $Y=80300 $D=8
D703 GND_PAD! VDD_PAD! dn PJ=0.00041 m=1 $X=7791540 $Y=80300 $D=8
D704 GND_PAD! VDD_PAD! dn PJ=0.00041 m=1 $X=7801540 $Y=80300 $D=8
D705 GND_PAD! VDD_PAD! dn PJ=0.00041 m=1 $X=7811540 $Y=80300 $D=8
D706 GND_PAD! VDD_PAD! dn PJ=0.00041 m=1 $X=7821540 $Y=80300 $D=8
D707 GND_PAD! VDD_PAD! dn PJ=0.00041 m=1 $X=7831540 $Y=80300 $D=8
D708 GND_PAD! VDD_PAD! dn PJ=0.00041 m=1 $X=7841540 $Y=80300 $D=8
D709 A13 vdd! dn PJ=0.0002 m=1 $X=10384020 $Y=13228100 $D=8
D710 A13 vdd! dn PJ=0.0002 m=1 $X=10384020 $Y=13438100 $D=8
D711 gnd! A13 dn PJ=0.0002 m=1 $X=10386340 $Y=13232500 $D=8
D712 gnd! A13 dn PJ=0.0002 m=1 $X=10386340 $Y=13442500 $D=8
D713 A13 vdd! dn PJ=0.0002 m=1 $X=10388660 $Y=13228100 $D=8
D714 A13 vdd! dn PJ=0.0002 m=1 $X=10388660 $Y=13438100 $D=8
D715 gnd! A13 dn PJ=0.0001 m=1 $X=10390980 $Y=13332500 $D=8
D716 gnd! A13 dn PJ=0.0001 m=1 $X=10390980 $Y=13542500 $D=8
D717 A13 vdd! dn PJ=0.0001 m=1 $X=10394160 $Y=13228100 $D=8
D718 A13 vdd! dn PJ=0.0001 m=1 $X=10394160 $Y=13438100 $D=8
D719 gnd! A13 dn PJ=0.0002 m=1 $X=10396480 $Y=13232500 $D=8
D720 gnd! A13 dn PJ=0.0002 m=1 $X=10396480 $Y=13442500 $D=8
D721 A13 vdd! dn PJ=0.0002 m=1 $X=10398800 $Y=13228100 $D=8
D722 A13 vdd! dn PJ=0.0002 m=1 $X=10398800 $Y=13438100 $D=8
D723 gnd! A13 dn PJ=0.0002 m=1 $X=10401120 $Y=13232500 $D=8
D724 gnd! A13 dn PJ=0.0002 m=1 $X=10401120 $Y=13442500 $D=8
D725 A13 vdd! dn PJ=0.0002 m=1 $X=10403440 $Y=13228100 $D=8
D726 A13 vdd! dn PJ=0.0002 m=1 $X=10403440 $Y=13438100 $D=8
D727 gnd! A13 dn PJ=0.0001 m=1 $X=10405760 $Y=13332500 $D=8
D728 gnd! A13 dn PJ=0.0001 m=1 $X=10405760 $Y=13542500 $D=8
D729 A13 vdd! dn PJ=0.0001 m=1 $X=10408940 $Y=13228100 $D=8
D730 A13 vdd! dn PJ=0.0001 m=1 $X=10408940 $Y=13438100 $D=8
D731 gnd! A13 dn PJ=0.0002 m=1 $X=10411260 $Y=13232500 $D=8
D732 gnd! A13 dn PJ=0.0002 m=1 $X=10411260 $Y=13442500 $D=8
D733 A13 vdd! dn PJ=0.0002 m=1 $X=10413580 $Y=13228100 $D=8
D734 A13 vdd! dn PJ=0.0002 m=1 $X=10413580 $Y=13438100 $D=8
D735 gnd! A13 dn PJ=0.0002 m=1 $X=10415900 $Y=13232500 $D=8
D736 gnd! A13 dn PJ=0.0002 m=1 $X=10415900 $Y=13442500 $D=8
D737 A13 vdd! dn PJ=0.0002 m=1 $X=10418220 $Y=13228100 $D=8
D738 A13 vdd! dn PJ=0.0002 m=1 $X=10418220 $Y=13438100 $D=8
D739 gnd! A13 dn PJ=0.0001 m=1 $X=10420540 $Y=13332500 $D=8
D740 gnd! A13 dn PJ=0.0001 m=1 $X=10420540 $Y=13542500 $D=8
D741 A13 vdd! dn PJ=0.0001 m=1 $X=10423720 $Y=13228100 $D=8
D742 A13 vdd! dn PJ=0.0001 m=1 $X=10423720 $Y=13438100 $D=8
D743 gnd! A13 dn PJ=0.0002 m=1 $X=10426040 $Y=13232500 $D=8
D744 gnd! A13 dn PJ=0.0002 m=1 $X=10426040 $Y=13442500 $D=8
D745 A13 vdd! dn PJ=0.0002 m=1 $X=10428360 $Y=13228100 $D=8
D746 A13 vdd! dn PJ=0.0002 m=1 $X=10428360 $Y=13438100 $D=8
D747 gnd! A13 dn PJ=0.0002 m=1 $X=10430680 $Y=13232500 $D=8
D748 gnd! A13 dn PJ=0.0002 m=1 $X=10430680 $Y=13442500 $D=8
D749 A13 vdd! dn PJ=0.0002 m=1 $X=10433000 $Y=13228100 $D=8
D750 A13 vdd! dn PJ=0.0002 m=1 $X=10433000 $Y=13438100 $D=8
D751 gnd! A13 dn PJ=0.0001 m=1 $X=10435320 $Y=13332500 $D=8
D752 gnd! A13 dn PJ=0.0001 m=1 $X=10435320 $Y=13542500 $D=8
D753 A13 vdd! dn PJ=0.0001 m=1 $X=10438500 $Y=13228100 $D=8
D754 A13 vdd! dn PJ=0.0001 m=1 $X=10438500 $Y=13438100 $D=8
D755 gnd! A13 dn PJ=0.0002 m=1 $X=10440820 $Y=13232500 $D=8
D756 gnd! A13 dn PJ=0.0002 m=1 $X=10440820 $Y=13442500 $D=8
D757 A13 vdd! dn PJ=0.0002 m=1 $X=10443140 $Y=13228100 $D=8
D758 A13 vdd! dn PJ=0.0002 m=1 $X=10443140 $Y=13438100 $D=8
D759 gnd! A13 dn PJ=0.0002 m=1 $X=10445460 $Y=13232500 $D=8
D760 gnd! A13 dn PJ=0.0002 m=1 $X=10445460 $Y=13442500 $D=8
D761 A13 vdd! dn PJ=0.0002 m=1 $X=10447780 $Y=13228100 $D=8
D762 A13 vdd! dn PJ=0.0002 m=1 $X=10447780 $Y=13438100 $D=8
D763 gnd! A13 dn PJ=0.0001 m=1 $X=10450100 $Y=13332500 $D=8
D764 gnd! A13 dn PJ=0.0001 m=1 $X=10450100 $Y=13542500 $D=8
D765 A13 vdd! dn PJ=0.0001 m=1 $X=10453280 $Y=13228100 $D=8
D766 A13 vdd! dn PJ=0.0001 m=1 $X=10453280 $Y=13438100 $D=8
D767 gnd! A13 dn PJ=0.0002 m=1 $X=10455600 $Y=13232500 $D=8
D768 gnd! A13 dn PJ=0.0002 m=1 $X=10455600 $Y=13442500 $D=8
D769 A13 vdd! dn PJ=0.0002 m=1 $X=10457920 $Y=13228100 $D=8
D770 A13 vdd! dn PJ=0.0002 m=1 $X=10457920 $Y=13438100 $D=8
D771 gnd! A13 dn PJ=0.0002 m=1 $X=10460240 $Y=13232500 $D=8
D772 gnd! A13 dn PJ=0.0002 m=1 $X=10460240 $Y=13442500 $D=8
D773 GND_PAD! VDD_PAD! dn PJ=0.00041 m=1 $X=10461540 $Y=80300 $D=8
D774 A13 vdd! dn PJ=0.0002 m=1 $X=10462560 $Y=13228100 $D=8
D775 A13 vdd! dn PJ=0.0002 m=1 $X=10462560 $Y=13438100 $D=8
D776 gnd! A13 dn PJ=0.0001 m=1 $X=10464880 $Y=13332500 $D=8
D777 gnd! A13 dn PJ=0.0001 m=1 $X=10464880 $Y=13542500 $D=8
D778 A13 vdd! dn PJ=0.0001 m=1 $X=10468060 $Y=13228100 $D=8
D779 A13 vdd! dn PJ=0.0001 m=1 $X=10468060 $Y=13438100 $D=8
D780 gnd! A13 dn PJ=0.0002 m=1 $X=10470380 $Y=13232500 $D=8
D781 gnd! A13 dn PJ=0.0002 m=1 $X=10470380 $Y=13442500 $D=8
D782 GND_PAD! VDD_PAD! dn PJ=0.00041 m=1 $X=10471540 $Y=80300 $D=8
D783 A13 vdd! dn PJ=0.0002 m=1 $X=10472700 $Y=13228100 $D=8
D784 A13 vdd! dn PJ=0.0002 m=1 $X=10472700 $Y=13438100 $D=8
D785 gnd! A13 dn PJ=0.0002 m=1 $X=10475020 $Y=13232500 $D=8
D786 gnd! A13 dn PJ=0.0002 m=1 $X=10475020 $Y=13442500 $D=8
D787 GND_PAD! VDD_PAD! dn PJ=0.00041 m=1 $X=10481540 $Y=80300 $D=8
D788 GND_PAD! VDD_PAD! dn PJ=0.00041 m=1 $X=10491540 $Y=80300 $D=8
D789 GND_PAD! VDD_PAD! dn PJ=0.00041 m=1 $X=10501540 $Y=80300 $D=8
D790 GND_PAD! VDD_PAD! dn PJ=0.00041 m=1 $X=10511540 $Y=80300 $D=8
D791 GND_PAD! VDD_PAD! dn PJ=0.00041 m=1 $X=10521540 $Y=80300 $D=8
D792 GND_PAD! VDD_PAD! dn PJ=0.00041 m=1 $X=10531540 $Y=80300 $D=8
D793 GND_PAD! VDD_PAD! dn PJ=0.00041 m=1 $X=10541540 $Y=80300 $D=8
D794 GND_PAD! VDD_PAD! dn PJ=0.00041 m=1 $X=10761540 $Y=80300 $D=8
D795 GND_PAD! VDD_PAD! dn PJ=0.00041 m=1 $X=10771540 $Y=80300 $D=8
D796 GND_PAD! VDD_PAD! dn PJ=0.00041 m=1 $X=10781540 $Y=80300 $D=8
D797 GND_PAD! VDD_PAD! dn PJ=0.00041 m=1 $X=10791540 $Y=80300 $D=8
D798 GND_PAD! VDD_PAD! dn PJ=0.00041 m=1 $X=10801540 $Y=80300 $D=8
D799 GND_PAD! VDD_PAD! dn PJ=0.00041 m=1 $X=10811540 $Y=80300 $D=8
D800 GND_PAD! VDD_PAD! dn PJ=0.00041 m=1 $X=10821540 $Y=80300 $D=8
D801 GND_PAD! VDD_PAD! dn PJ=0.00041 m=1 $X=10831540 $Y=80300 $D=8
D802 GND_PAD! VDD_PAD! dn PJ=0.00041 m=1 $X=10841540 $Y=80300 $D=8
D803 A15 vdd! dn PJ=0.0002 m=1 $X=10904020 $Y=13228100 $D=8
D804 A15 vdd! dn PJ=0.0002 m=1 $X=10904020 $Y=13438100 $D=8
D805 gnd! A15 dn PJ=0.0002 m=1 $X=10906340 $Y=13232500 $D=8
D806 gnd! A15 dn PJ=0.0002 m=1 $X=10906340 $Y=13442500 $D=8
D807 A15 vdd! dn PJ=0.0002 m=1 $X=10908660 $Y=13228100 $D=8
D808 A15 vdd! dn PJ=0.0002 m=1 $X=10908660 $Y=13438100 $D=8
D809 gnd! A15 dn PJ=0.0001 m=1 $X=10910980 $Y=13332500 $D=8
D810 gnd! A15 dn PJ=0.0001 m=1 $X=10910980 $Y=13542500 $D=8
D811 A15 vdd! dn PJ=0.0001 m=1 $X=10914160 $Y=13228100 $D=8
D812 A15 vdd! dn PJ=0.0001 m=1 $X=10914160 $Y=13438100 $D=8
D813 gnd! A15 dn PJ=0.0002 m=1 $X=10916480 $Y=13232500 $D=8
D814 gnd! A15 dn PJ=0.0002 m=1 $X=10916480 $Y=13442500 $D=8
D815 A15 vdd! dn PJ=0.0002 m=1 $X=10918800 $Y=13228100 $D=8
D816 A15 vdd! dn PJ=0.0002 m=1 $X=10918800 $Y=13438100 $D=8
D817 gnd! A15 dn PJ=0.0002 m=1 $X=10921120 $Y=13232500 $D=8
D818 gnd! A15 dn PJ=0.0002 m=1 $X=10921120 $Y=13442500 $D=8
D819 A15 vdd! dn PJ=0.0002 m=1 $X=10923440 $Y=13228100 $D=8
D820 A15 vdd! dn PJ=0.0002 m=1 $X=10923440 $Y=13438100 $D=8
D821 gnd! A15 dn PJ=0.0001 m=1 $X=10925760 $Y=13332500 $D=8
D822 gnd! A15 dn PJ=0.0001 m=1 $X=10925760 $Y=13542500 $D=8
D823 A15 vdd! dn PJ=0.0001 m=1 $X=10928940 $Y=13228100 $D=8
D824 A15 vdd! dn PJ=0.0001 m=1 $X=10928940 $Y=13438100 $D=8
D825 gnd! A15 dn PJ=0.0002 m=1 $X=10931260 $Y=13232500 $D=8
D826 gnd! A15 dn PJ=0.0002 m=1 $X=10931260 $Y=13442500 $D=8
D827 A15 vdd! dn PJ=0.0002 m=1 $X=10933580 $Y=13228100 $D=8
D828 A15 vdd! dn PJ=0.0002 m=1 $X=10933580 $Y=13438100 $D=8
D829 gnd! A15 dn PJ=0.0002 m=1 $X=10935900 $Y=13232500 $D=8
D830 gnd! A15 dn PJ=0.0002 m=1 $X=10935900 $Y=13442500 $D=8
D831 A15 vdd! dn PJ=0.0002 m=1 $X=10938220 $Y=13228100 $D=8
D832 A15 vdd! dn PJ=0.0002 m=1 $X=10938220 $Y=13438100 $D=8
D833 gnd! A15 dn PJ=0.0001 m=1 $X=10940540 $Y=13332500 $D=8
D834 gnd! A15 dn PJ=0.0001 m=1 $X=10940540 $Y=13542500 $D=8
D835 A15 vdd! dn PJ=0.0001 m=1 $X=10943720 $Y=13228100 $D=8
D836 A15 vdd! dn PJ=0.0001 m=1 $X=10943720 $Y=13438100 $D=8
D837 gnd! A15 dn PJ=0.0002 m=1 $X=10946040 $Y=13232500 $D=8
D838 gnd! A15 dn PJ=0.0002 m=1 $X=10946040 $Y=13442500 $D=8
D839 A15 vdd! dn PJ=0.0002 m=1 $X=10948360 $Y=13228100 $D=8
D840 A15 vdd! dn PJ=0.0002 m=1 $X=10948360 $Y=13438100 $D=8
D841 gnd! A15 dn PJ=0.0002 m=1 $X=10950680 $Y=13232500 $D=8
D842 gnd! A15 dn PJ=0.0002 m=1 $X=10950680 $Y=13442500 $D=8
D843 A15 vdd! dn PJ=0.0002 m=1 $X=10953000 $Y=13228100 $D=8
D844 A15 vdd! dn PJ=0.0002 m=1 $X=10953000 $Y=13438100 $D=8
D845 gnd! A15 dn PJ=0.0001 m=1 $X=10955320 $Y=13332500 $D=8
D846 gnd! A15 dn PJ=0.0001 m=1 $X=10955320 $Y=13542500 $D=8
D847 A15 vdd! dn PJ=0.0001 m=1 $X=10958500 $Y=13228100 $D=8
D848 A15 vdd! dn PJ=0.0001 m=1 $X=10958500 $Y=13438100 $D=8
D849 gnd! A15 dn PJ=0.0002 m=1 $X=10960820 $Y=13232500 $D=8
D850 gnd! A15 dn PJ=0.0002 m=1 $X=10960820 $Y=13442500 $D=8
D851 A15 vdd! dn PJ=0.0002 m=1 $X=10963140 $Y=13228100 $D=8
D852 A15 vdd! dn PJ=0.0002 m=1 $X=10963140 $Y=13438100 $D=8
D853 gnd! A15 dn PJ=0.0002 m=1 $X=10965460 $Y=13232500 $D=8
D854 gnd! A15 dn PJ=0.0002 m=1 $X=10965460 $Y=13442500 $D=8
D855 A15 vdd! dn PJ=0.0002 m=1 $X=10967780 $Y=13228100 $D=8
D856 A15 vdd! dn PJ=0.0002 m=1 $X=10967780 $Y=13438100 $D=8
D857 gnd! A15 dn PJ=0.0001 m=1 $X=10970100 $Y=13332500 $D=8
D858 gnd! A15 dn PJ=0.0001 m=1 $X=10970100 $Y=13542500 $D=8
D859 A15 vdd! dn PJ=0.0001 m=1 $X=10973280 $Y=13228100 $D=8
D860 A15 vdd! dn PJ=0.0001 m=1 $X=10973280 $Y=13438100 $D=8
D861 gnd! A15 dn PJ=0.0002 m=1 $X=10975600 $Y=13232500 $D=8
D862 gnd! A15 dn PJ=0.0002 m=1 $X=10975600 $Y=13442500 $D=8
D863 A15 vdd! dn PJ=0.0002 m=1 $X=10977920 $Y=13228100 $D=8
D864 A15 vdd! dn PJ=0.0002 m=1 $X=10977920 $Y=13438100 $D=8
D865 gnd! A15 dn PJ=0.0002 m=1 $X=10980240 $Y=13232500 $D=8
D866 gnd! A15 dn PJ=0.0002 m=1 $X=10980240 $Y=13442500 $D=8
D867 A15 vdd! dn PJ=0.0002 m=1 $X=10982560 $Y=13228100 $D=8
D868 A15 vdd! dn PJ=0.0002 m=1 $X=10982560 $Y=13438100 $D=8
D869 gnd! A15 dn PJ=0.0001 m=1 $X=10984880 $Y=13332500 $D=8
D870 gnd! A15 dn PJ=0.0001 m=1 $X=10984880 $Y=13542500 $D=8
D871 A15 vdd! dn PJ=0.0001 m=1 $X=10988060 $Y=13228100 $D=8
D872 A15 vdd! dn PJ=0.0001 m=1 $X=10988060 $Y=13438100 $D=8
D873 gnd! A15 dn PJ=0.0002 m=1 $X=10990380 $Y=13232500 $D=8
D874 gnd! A15 dn PJ=0.0002 m=1 $X=10990380 $Y=13442500 $D=8
D875 A15 vdd! dn PJ=0.0002 m=1 $X=10992700 $Y=13228100 $D=8
D876 A15 vdd! dn PJ=0.0002 m=1 $X=10992700 $Y=13438100 $D=8
D877 gnd! A15 dn PJ=0.0002 m=1 $X=10995020 $Y=13232500 $D=8
D878 gnd! A15 dn PJ=0.0002 m=1 $X=10995020 $Y=13442500 $D=8
D879 A16 vdd! dn PJ=0.0002 m=1 $X=11684020 $Y=13228100 $D=8
D880 A16 vdd! dn PJ=0.0002 m=1 $X=11684020 $Y=13438100 $D=8
D881 gnd! A16 dn PJ=0.0002 m=1 $X=11686340 $Y=13232500 $D=8
D882 gnd! A16 dn PJ=0.0002 m=1 $X=11686340 $Y=13442500 $D=8
D883 A16 vdd! dn PJ=0.0002 m=1 $X=11688660 $Y=13228100 $D=8
D884 A16 vdd! dn PJ=0.0002 m=1 $X=11688660 $Y=13438100 $D=8
D885 gnd! A16 dn PJ=0.0001 m=1 $X=11690980 $Y=13332500 $D=8
D886 gnd! A16 dn PJ=0.0001 m=1 $X=11690980 $Y=13542500 $D=8
D887 A16 vdd! dn PJ=0.0001 m=1 $X=11694160 $Y=13228100 $D=8
D888 A16 vdd! dn PJ=0.0001 m=1 $X=11694160 $Y=13438100 $D=8
D889 gnd! A16 dn PJ=0.0002 m=1 $X=11696480 $Y=13232500 $D=8
D890 gnd! A16 dn PJ=0.0002 m=1 $X=11696480 $Y=13442500 $D=8
D891 A16 vdd! dn PJ=0.0002 m=1 $X=11698800 $Y=13228100 $D=8
D892 A16 vdd! dn PJ=0.0002 m=1 $X=11698800 $Y=13438100 $D=8
D893 gnd! A16 dn PJ=0.0002 m=1 $X=11701120 $Y=13232500 $D=8
D894 gnd! A16 dn PJ=0.0002 m=1 $X=11701120 $Y=13442500 $D=8
D895 A16 vdd! dn PJ=0.0002 m=1 $X=11703440 $Y=13228100 $D=8
D896 A16 vdd! dn PJ=0.0002 m=1 $X=11703440 $Y=13438100 $D=8
D897 gnd! A16 dn PJ=0.0001 m=1 $X=11705760 $Y=13332500 $D=8
D898 gnd! A16 dn PJ=0.0001 m=1 $X=11705760 $Y=13542500 $D=8
D899 A16 vdd! dn PJ=0.0001 m=1 $X=11708940 $Y=13228100 $D=8
D900 A16 vdd! dn PJ=0.0001 m=1 $X=11708940 $Y=13438100 $D=8
D901 gnd! A16 dn PJ=0.0002 m=1 $X=11711260 $Y=13232500 $D=8
D902 gnd! A16 dn PJ=0.0002 m=1 $X=11711260 $Y=13442500 $D=8
D903 A16 vdd! dn PJ=0.0002 m=1 $X=11713580 $Y=13228100 $D=8
D904 A16 vdd! dn PJ=0.0002 m=1 $X=11713580 $Y=13438100 $D=8
D905 gnd! A16 dn PJ=0.0002 m=1 $X=11715900 $Y=13232500 $D=8
D906 gnd! A16 dn PJ=0.0002 m=1 $X=11715900 $Y=13442500 $D=8
D907 A16 vdd! dn PJ=0.0002 m=1 $X=11718220 $Y=13228100 $D=8
D908 A16 vdd! dn PJ=0.0002 m=1 $X=11718220 $Y=13438100 $D=8
D909 gnd! A16 dn PJ=0.0001 m=1 $X=11720540 $Y=13332500 $D=8
D910 gnd! A16 dn PJ=0.0001 m=1 $X=11720540 $Y=13542500 $D=8
D911 A16 vdd! dn PJ=0.0001 m=1 $X=11723720 $Y=13228100 $D=8
D912 A16 vdd! dn PJ=0.0001 m=1 $X=11723720 $Y=13438100 $D=8
D913 gnd! A16 dn PJ=0.0002 m=1 $X=11726040 $Y=13232500 $D=8
D914 gnd! A16 dn PJ=0.0002 m=1 $X=11726040 $Y=13442500 $D=8
D915 A16 vdd! dn PJ=0.0002 m=1 $X=11728360 $Y=13228100 $D=8
D916 A16 vdd! dn PJ=0.0002 m=1 $X=11728360 $Y=13438100 $D=8
D917 gnd! A16 dn PJ=0.0002 m=1 $X=11730680 $Y=13232500 $D=8
D918 gnd! A16 dn PJ=0.0002 m=1 $X=11730680 $Y=13442500 $D=8
D919 A16 vdd! dn PJ=0.0002 m=1 $X=11733000 $Y=13228100 $D=8
D920 A16 vdd! dn PJ=0.0002 m=1 $X=11733000 $Y=13438100 $D=8
D921 gnd! A16 dn PJ=0.0001 m=1 $X=11735320 $Y=13332500 $D=8
D922 gnd! A16 dn PJ=0.0001 m=1 $X=11735320 $Y=13542500 $D=8
D923 A16 vdd! dn PJ=0.0001 m=1 $X=11738500 $Y=13228100 $D=8
D924 A16 vdd! dn PJ=0.0001 m=1 $X=11738500 $Y=13438100 $D=8
D925 gnd! A16 dn PJ=0.0002 m=1 $X=11740820 $Y=13232500 $D=8
D926 gnd! A16 dn PJ=0.0002 m=1 $X=11740820 $Y=13442500 $D=8
D927 A16 vdd! dn PJ=0.0002 m=1 $X=11743140 $Y=13228100 $D=8
D928 A16 vdd! dn PJ=0.0002 m=1 $X=11743140 $Y=13438100 $D=8
D929 gnd! A16 dn PJ=0.0002 m=1 $X=11745460 $Y=13232500 $D=8
D930 gnd! A16 dn PJ=0.0002 m=1 $X=11745460 $Y=13442500 $D=8
D931 A16 vdd! dn PJ=0.0002 m=1 $X=11747780 $Y=13228100 $D=8
D932 A16 vdd! dn PJ=0.0002 m=1 $X=11747780 $Y=13438100 $D=8
D933 gnd! A16 dn PJ=0.0001 m=1 $X=11750100 $Y=13332500 $D=8
D934 gnd! A16 dn PJ=0.0001 m=1 $X=11750100 $Y=13542500 $D=8
D935 A16 vdd! dn PJ=0.0001 m=1 $X=11753280 $Y=13228100 $D=8
D936 A16 vdd! dn PJ=0.0001 m=1 $X=11753280 $Y=13438100 $D=8
D937 gnd! A16 dn PJ=0.0002 m=1 $X=11755600 $Y=13232500 $D=8
D938 gnd! A16 dn PJ=0.0002 m=1 $X=11755600 $Y=13442500 $D=8
D939 A16 vdd! dn PJ=0.0002 m=1 $X=11757920 $Y=13228100 $D=8
D940 A16 vdd! dn PJ=0.0002 m=1 $X=11757920 $Y=13438100 $D=8
D941 gnd! A16 dn PJ=0.0002 m=1 $X=11760240 $Y=13232500 $D=8
D942 gnd! A16 dn PJ=0.0002 m=1 $X=11760240 $Y=13442500 $D=8
D943 A16 vdd! dn PJ=0.0002 m=1 $X=11762560 $Y=13228100 $D=8
D944 A16 vdd! dn PJ=0.0002 m=1 $X=11762560 $Y=13438100 $D=8
D945 gnd! A16 dn PJ=0.0001 m=1 $X=11764880 $Y=13332500 $D=8
D946 gnd! A16 dn PJ=0.0001 m=1 $X=11764880 $Y=13542500 $D=8
D947 A16 vdd! dn PJ=0.0001 m=1 $X=11768060 $Y=13228100 $D=8
D948 A16 vdd! dn PJ=0.0001 m=1 $X=11768060 $Y=13438100 $D=8
D949 gnd! A16 dn PJ=0.0002 m=1 $X=11770380 $Y=13232500 $D=8
D950 gnd! A16 dn PJ=0.0002 m=1 $X=11770380 $Y=13442500 $D=8
D951 A16 vdd! dn PJ=0.0002 m=1 $X=11772700 $Y=13228100 $D=8
D952 A16 vdd! dn PJ=0.0002 m=1 $X=11772700 $Y=13438100 $D=8
D953 gnd! A16 dn PJ=0.0002 m=1 $X=11775020 $Y=13232500 $D=8
D954 gnd! A16 dn PJ=0.0002 m=1 $X=11775020 $Y=13442500 $D=8
D955 GND_PAD! VDD_PAD! dn PJ=0.00041 m=1 $X=14061540 $Y=80300 $D=8
D956 GND_PAD! VDD_PAD! dn PJ=0.00041 m=1 $X=14071540 $Y=80300 $D=8
D957 GND_PAD! VDD_PAD! dn PJ=0.00041 m=1 $X=14081540 $Y=80300 $D=8
D958 GND_PAD! VDD_PAD! dn PJ=0.00041 m=1 $X=14091540 $Y=80300 $D=8
D959 GND_PAD! VDD_PAD! dn PJ=0.00041 m=1 $X=14101540 $Y=80300 $D=8
D960 GND_PAD! VDD_PAD! dn PJ=0.00041 m=1 $X=14111540 $Y=80300 $D=8
D961 GND_PAD! VDD_PAD! dn PJ=0.00041 m=1 $X=14121540 $Y=80300 $D=8
D962 GND_PAD! VDD_PAD! dn PJ=0.00041 m=1 $X=14131540 $Y=80300 $D=8
D963 GND_PAD! VDD_PAD! dn PJ=0.00041 m=1 $X=14141540 $Y=80300 $D=8
D964 GND_PAD! VDD_PAD! dn PJ=0.00041 m=1 $X=-45240 $Y=80300 $D=9
D965 VDD_PAD! vdd! dn PJ=0.00041 m=1 $X=-42740 $Y=80300 $D=9
D966 vdd! VDD_PAD! dn PJ=0.00041 m=1 $X=-40240 $Y=80300 $D=9
D967 GND_PAD! VDD_PAD! dn PJ=0.00041 m=1 $X=-35240 $Y=80300 $D=9
D968 VDD_PAD! vdd! dn PJ=0.00041 m=1 $X=-32740 $Y=80300 $D=9
D969 vdd! VDD_PAD! dn PJ=0.00041 m=1 $X=-30240 $Y=80300 $D=9
D970 GND_PAD! VDD_PAD! dn PJ=0.00041 m=1 $X=-25240 $Y=80300 $D=9
D971 VDD_PAD! vdd! dn PJ=0.00041 m=1 $X=-22740 $Y=80300 $D=9
D972 vdd! VDD_PAD! dn PJ=0.00041 m=1 $X=-20240 $Y=80300 $D=9
D973 gnd! Test dn PJ=0.0002 m=1 $X=-16000 $Y=13232500 $D=9
D974 gnd! Test dn PJ=0.0002 m=1 $X=-16000 $Y=13442500 $D=9
D975 GND_PAD! VDD_PAD! dn PJ=0.00041 m=1 $X=-15240 $Y=80300 $D=9
D976 Test vdd! dn PJ=0.0002 m=1 $X=-13680 $Y=13228100 $D=9
D977 Test vdd! dn PJ=0.0002 m=1 $X=-13680 $Y=13438100 $D=9
D978 VDD_PAD! vdd! dn PJ=0.00041 m=1 $X=-12740 $Y=80300 $D=9
D979 gnd! Test dn PJ=0.0002 m=1 $X=-11360 $Y=13232500 $D=9
D980 gnd! Test dn PJ=0.0002 m=1 $X=-11360 $Y=13442500 $D=9
D981 vdd! VDD_PAD! dn PJ=0.00041 m=1 $X=-10240 $Y=80300 $D=9
D982 Test vdd! dn PJ=0.0001 m=1 $X=-9040 $Y=13228100 $D=9
D983 Test vdd! dn PJ=0.0001 m=1 $X=-9040 $Y=13438100 $D=9
D984 gnd! Test dn PJ=0.0001 m=1 $X=-5860 $Y=13332500 $D=9
D985 gnd! Test dn PJ=0.0001 m=1 $X=-5860 $Y=13542500 $D=9
D986 GND_PAD! VDD_PAD! dn PJ=0.00041 m=1 $X=-5240 $Y=80300 $D=9
D987 Test vdd! dn PJ=0.0002 m=1 $X=-3540 $Y=13228100 $D=9
D988 Test vdd! dn PJ=0.0002 m=1 $X=-3540 $Y=13438100 $D=9
D989 VDD_PAD! vdd! dn PJ=0.00041 m=1 $X=-2740 $Y=80300 $D=9
D990 gnd! Test dn PJ=0.0002 m=1 $X=-1220 $Y=13232500 $D=9
D991 gnd! Test dn PJ=0.0002 m=1 $X=-1220 $Y=13442500 $D=9
D992 vdd! VDD_PAD! dn PJ=0.00041 m=1 $X=-240 $Y=80300 $D=9
D993 Test vdd! dn PJ=0.0002 m=1 $X=1100 $Y=13228100 $D=9
D994 Test vdd! dn PJ=0.0002 m=1 $X=1100 $Y=13438100 $D=9
D995 gnd! Test dn PJ=0.0002 m=1 $X=3420 $Y=13232500 $D=9
D996 gnd! Test dn PJ=0.0002 m=1 $X=3420 $Y=13442500 $D=9
D997 GND_PAD! VDD_PAD! dn PJ=0.00041 m=1 $X=4760 $Y=80300 $D=9
D998 Test vdd! dn PJ=0.0001 m=1 $X=5740 $Y=13228100 $D=9
D999 Test vdd! dn PJ=0.0001 m=1 $X=5740 $Y=13438100 $D=9
D1000 VDD_PAD! vdd! dn PJ=0.00041 m=1 $X=7260 $Y=80300 $D=9
D1001 gnd! Test dn PJ=0.0001 m=1 $X=8920 $Y=13332500 $D=9
D1002 gnd! Test dn PJ=0.0001 m=1 $X=8920 $Y=13542500 $D=9
D1003 vdd! VDD_PAD! dn PJ=0.00041 m=1 $X=9760 $Y=80300 $D=9
D1004 Test vdd! dn PJ=0.0002 m=1 $X=11240 $Y=13228100 $D=9
D1005 Test vdd! dn PJ=0.0002 m=1 $X=11240 $Y=13438100 $D=9
D1006 gnd! Test dn PJ=0.0002 m=1 $X=13560 $Y=13232500 $D=9
D1007 gnd! Test dn PJ=0.0002 m=1 $X=13560 $Y=13442500 $D=9
D1008 GND_PAD! VDD_PAD! dn PJ=0.00041 m=1 $X=14760 $Y=80300 $D=9
D1009 Test vdd! dn PJ=0.0002 m=1 $X=15880 $Y=13228100 $D=9
D1010 Test vdd! dn PJ=0.0002 m=1 $X=15880 $Y=13438100 $D=9
D1011 VDD_PAD! vdd! dn PJ=0.00041 m=1 $X=17260 $Y=80300 $D=9
D1012 gnd! Test dn PJ=0.0002 m=1 $X=18200 $Y=13232500 $D=9
D1013 gnd! Test dn PJ=0.0002 m=1 $X=18200 $Y=13442500 $D=9
D1014 vdd! VDD_PAD! dn PJ=0.00041 m=1 $X=19760 $Y=80300 $D=9
D1015 Test vdd! dn PJ=0.0001 m=1 $X=20520 $Y=13228100 $D=9
D1016 Test vdd! dn PJ=0.0001 m=1 $X=20520 $Y=13438100 $D=9
D1017 gnd! Test dn PJ=0.0001 m=1 $X=23700 $Y=13332500 $D=9
D1018 gnd! Test dn PJ=0.0001 m=1 $X=23700 $Y=13542500 $D=9
D1019 GND_PAD! VDD_PAD! dn PJ=0.00041 m=1 $X=24760 $Y=80300 $D=9
D1020 Test vdd! dn PJ=0.0002 m=1 $X=26020 $Y=13228100 $D=9
D1021 Test vdd! dn PJ=0.0002 m=1 $X=26020 $Y=13438100 $D=9
D1022 VDD_PAD! vdd! dn PJ=0.00041 m=1 $X=27260 $Y=80300 $D=9
D1023 gnd! Test dn PJ=0.0002 m=1 $X=28340 $Y=13232500 $D=9
D1024 gnd! Test dn PJ=0.0002 m=1 $X=28340 $Y=13442500 $D=9
D1025 vdd! VDD_PAD! dn PJ=0.00041 m=1 $X=29760 $Y=80300 $D=9
D1026 Test vdd! dn PJ=0.0002 m=1 $X=30660 $Y=13228100 $D=9
D1027 Test vdd! dn PJ=0.0002 m=1 $X=30660 $Y=13438100 $D=9
D1028 gnd! Test dn PJ=0.0002 m=1 $X=32980 $Y=13232500 $D=9
D1029 gnd! Test dn PJ=0.0002 m=1 $X=32980 $Y=13442500 $D=9
D1030 GND_PAD! VDD_PAD! dn PJ=0.00041 m=1 $X=34760 $Y=80300 $D=9
D1031 Test vdd! dn PJ=0.0001 m=1 $X=35300 $Y=13228100 $D=9
D1032 Test vdd! dn PJ=0.0001 m=1 $X=35300 $Y=13438100 $D=9
D1033 VDD_PAD! vdd! dn PJ=0.00041 m=1 $X=37260 $Y=80300 $D=9
D1034 gnd! Test dn PJ=0.0001 m=1 $X=38480 $Y=13332500 $D=9
D1035 gnd! Test dn PJ=0.0001 m=1 $X=38480 $Y=13542500 $D=9
D1036 vdd! VDD_PAD! dn PJ=0.00041 m=1 $X=39760 $Y=80300 $D=9
D1037 Test vdd! dn PJ=0.0002 m=1 $X=40800 $Y=13228100 $D=9
D1038 Test vdd! dn PJ=0.0002 m=1 $X=40800 $Y=13438100 $D=9
D1039 gnd! Test dn PJ=0.0002 m=1 $X=43120 $Y=13232500 $D=9
D1040 gnd! Test dn PJ=0.0002 m=1 $X=43120 $Y=13442500 $D=9
D1041 GND_PAD! VDD_PAD! dn PJ=0.00041 m=1 $X=44760 $Y=80300 $D=9
D1042 Test vdd! dn PJ=0.0002 m=1 $X=45440 $Y=13228100 $D=9
D1043 Test vdd! dn PJ=0.0002 m=1 $X=45440 $Y=13438100 $D=9
D1044 VDD_PAD! vdd! dn PJ=0.00041 m=1 $X=47260 $Y=80300 $D=9
D1045 gnd! Test dn PJ=0.0002 m=1 $X=47760 $Y=13232500 $D=9
D1046 gnd! Test dn PJ=0.0002 m=1 $X=47760 $Y=13442500 $D=9
D1047 Test vdd! dn PJ=0.0001 m=1 $X=50080 $Y=13228100 $D=9
D1048 Test vdd! dn PJ=0.0001 m=1 $X=50080 $Y=13438100 $D=9
D1049 gnd! Test dn PJ=0.0001 m=1 $X=53260 $Y=13332500 $D=9
D1050 gnd! Test dn PJ=0.0001 m=1 $X=53260 $Y=13542500 $D=9
D1051 Test vdd! dn PJ=0.0002 m=1 $X=55580 $Y=13228100 $D=9
D1052 Test vdd! dn PJ=0.0002 m=1 $X=55580 $Y=13438100 $D=9
D1053 gnd! Test dn PJ=0.0002 m=1 $X=57900 $Y=13232500 $D=9
D1054 gnd! Test dn PJ=0.0002 m=1 $X=57900 $Y=13442500 $D=9
D1055 Test vdd! dn PJ=0.0002 m=1 $X=60220 $Y=13228100 $D=9
D1056 Test vdd! dn PJ=0.0002 m=1 $X=60220 $Y=13438100 $D=9
D1057 gnd! Test dn PJ=0.0002 m=1 $X=62540 $Y=13232500 $D=9
D1058 gnd! Test dn PJ=0.0002 m=1 $X=62540 $Y=13442500 $D=9
D1059 Test vdd! dn PJ=0.0001 m=1 $X=64860 $Y=13228100 $D=9
D1060 Test vdd! dn PJ=0.0001 m=1 $X=64860 $Y=13438100 $D=9
D1061 gnd! Test dn PJ=0.0001 m=1 $X=68040 $Y=13332500 $D=9
D1062 gnd! Test dn PJ=0.0001 m=1 $X=68040 $Y=13542500 $D=9
D1063 Test vdd! dn PJ=0.0002 m=1 $X=70360 $Y=13228100 $D=9
D1064 Test vdd! dn PJ=0.0002 m=1 $X=70360 $Y=13438100 $D=9
D1065 gnd! Test dn PJ=0.0002 m=1 $X=72680 $Y=13232500 $D=9
D1066 gnd! Test dn PJ=0.0002 m=1 $X=72680 $Y=13442500 $D=9
D1067 Test vdd! dn PJ=0.0002 m=1 $X=75000 $Y=13228100 $D=9
D1068 Test vdd! dn PJ=0.0002 m=1 $X=75000 $Y=13438100 $D=9
D1069 gnd! 252 dn PJ=0.0002 m=1 $X=244000 $Y=13232500 $D=9
D1070 gnd! 252 dn PJ=0.0002 m=1 $X=244000 $Y=13442500 $D=9
D1071 252 vdd! dn PJ=0.0002 m=1 $X=246320 $Y=13228100 $D=9
D1072 252 vdd! dn PJ=0.0002 m=1 $X=246320 $Y=13438100 $D=9
D1073 gnd! 252 dn PJ=0.0002 m=1 $X=248640 $Y=13232500 $D=9
D1074 gnd! 252 dn PJ=0.0002 m=1 $X=248640 $Y=13442500 $D=9
D1075 252 vdd! dn PJ=0.0001 m=1 $X=250960 $Y=13228100 $D=9
D1076 252 vdd! dn PJ=0.0001 m=1 $X=250960 $Y=13438100 $D=9
D1077 gnd! 252 dn PJ=0.0001 m=1 $X=254140 $Y=13332500 $D=9
D1078 gnd! 252 dn PJ=0.0001 m=1 $X=254140 $Y=13542500 $D=9
D1079 252 vdd! dn PJ=0.0002 m=1 $X=256460 $Y=13228100 $D=9
D1080 252 vdd! dn PJ=0.0002 m=1 $X=256460 $Y=13438100 $D=9
D1081 gnd! 252 dn PJ=0.0002 m=1 $X=258780 $Y=13232500 $D=9
D1082 gnd! 252 dn PJ=0.0002 m=1 $X=258780 $Y=13442500 $D=9
D1083 252 vdd! dn PJ=0.0002 m=1 $X=261100 $Y=13228100 $D=9
D1084 252 vdd! dn PJ=0.0002 m=1 $X=261100 $Y=13438100 $D=9
D1085 gnd! 252 dn PJ=0.0002 m=1 $X=263420 $Y=13232500 $D=9
D1086 gnd! 252 dn PJ=0.0002 m=1 $X=263420 $Y=13442500 $D=9
D1087 252 vdd! dn PJ=0.0001 m=1 $X=265740 $Y=13228100 $D=9
D1088 252 vdd! dn PJ=0.0001 m=1 $X=265740 $Y=13438100 $D=9
D1089 gnd! 252 dn PJ=0.0001 m=1 $X=268920 $Y=13332500 $D=9
D1090 gnd! 252 dn PJ=0.0001 m=1 $X=268920 $Y=13542500 $D=9
D1091 252 vdd! dn PJ=0.0002 m=1 $X=271240 $Y=13228100 $D=9
D1092 252 vdd! dn PJ=0.0002 m=1 $X=271240 $Y=13438100 $D=9
D1093 gnd! 252 dn PJ=0.0002 m=1 $X=273560 $Y=13232500 $D=9
D1094 gnd! 252 dn PJ=0.0002 m=1 $X=273560 $Y=13442500 $D=9
D1095 252 vdd! dn PJ=0.0002 m=1 $X=275880 $Y=13228100 $D=9
D1096 252 vdd! dn PJ=0.0002 m=1 $X=275880 $Y=13438100 $D=9
D1097 gnd! 252 dn PJ=0.0002 m=1 $X=278200 $Y=13232500 $D=9
D1098 gnd! 252 dn PJ=0.0002 m=1 $X=278200 $Y=13442500 $D=9
D1099 252 vdd! dn PJ=0.0001 m=1 $X=280520 $Y=13228100 $D=9
D1100 252 vdd! dn PJ=0.0001 m=1 $X=280520 $Y=13438100 $D=9
D1101 gnd! 252 dn PJ=0.0001 m=1 $X=283700 $Y=13332500 $D=9
D1102 gnd! 252 dn PJ=0.0001 m=1 $X=283700 $Y=13542500 $D=9
D1103 252 vdd! dn PJ=0.0002 m=1 $X=286020 $Y=13228100 $D=9
D1104 252 vdd! dn PJ=0.0002 m=1 $X=286020 $Y=13438100 $D=9
D1105 gnd! 252 dn PJ=0.0002 m=1 $X=288340 $Y=13232500 $D=9
D1106 gnd! 252 dn PJ=0.0002 m=1 $X=288340 $Y=13442500 $D=9
D1107 252 vdd! dn PJ=0.0002 m=1 $X=290660 $Y=13228100 $D=9
D1108 252 vdd! dn PJ=0.0002 m=1 $X=290660 $Y=13438100 $D=9
D1109 gnd! 252 dn PJ=0.0002 m=1 $X=292980 $Y=13232500 $D=9
D1110 gnd! 252 dn PJ=0.0002 m=1 $X=292980 $Y=13442500 $D=9
D1111 252 vdd! dn PJ=0.0001 m=1 $X=295300 $Y=13228100 $D=9
D1112 252 vdd! dn PJ=0.0001 m=1 $X=295300 $Y=13438100 $D=9
D1113 gnd! 252 dn PJ=0.0001 m=1 $X=298480 $Y=13332500 $D=9
D1114 gnd! 252 dn PJ=0.0001 m=1 $X=298480 $Y=13542500 $D=9
D1115 252 vdd! dn PJ=0.0002 m=1 $X=300800 $Y=13228100 $D=9
D1116 252 vdd! dn PJ=0.0002 m=1 $X=300800 $Y=13438100 $D=9
D1117 gnd! 252 dn PJ=0.0002 m=1 $X=303120 $Y=13232500 $D=9
D1118 gnd! 252 dn PJ=0.0002 m=1 $X=303120 $Y=13442500 $D=9
D1119 252 vdd! dn PJ=0.0002 m=1 $X=305440 $Y=13228100 $D=9
D1120 252 vdd! dn PJ=0.0002 m=1 $X=305440 $Y=13438100 $D=9
D1121 gnd! 252 dn PJ=0.0002 m=1 $X=307760 $Y=13232500 $D=9
D1122 gnd! 252 dn PJ=0.0002 m=1 $X=307760 $Y=13442500 $D=9
D1123 252 vdd! dn PJ=0.0001 m=1 $X=310080 $Y=13228100 $D=9
D1124 252 vdd! dn PJ=0.0001 m=1 $X=310080 $Y=13438100 $D=9
D1125 gnd! 252 dn PJ=0.0001 m=1 $X=313260 $Y=13332500 $D=9
D1126 gnd! 252 dn PJ=0.0001 m=1 $X=313260 $Y=13542500 $D=9
D1127 252 vdd! dn PJ=0.0002 m=1 $X=315580 $Y=13228100 $D=9
D1128 252 vdd! dn PJ=0.0002 m=1 $X=315580 $Y=13438100 $D=9
D1129 gnd! 252 dn PJ=0.0002 m=1 $X=317900 $Y=13232500 $D=9
D1130 gnd! 252 dn PJ=0.0002 m=1 $X=317900 $Y=13442500 $D=9
D1131 252 vdd! dn PJ=0.0002 m=1 $X=320220 $Y=13228100 $D=9
D1132 252 vdd! dn PJ=0.0002 m=1 $X=320220 $Y=13438100 $D=9
D1133 gnd! 252 dn PJ=0.0002 m=1 $X=322540 $Y=13232500 $D=9
D1134 gnd! 252 dn PJ=0.0002 m=1 $X=322540 $Y=13442500 $D=9
D1135 252 vdd! dn PJ=0.0001 m=1 $X=324860 $Y=13228100 $D=9
D1136 252 vdd! dn PJ=0.0001 m=1 $X=324860 $Y=13438100 $D=9
D1137 gnd! 252 dn PJ=0.0001 m=1 $X=328040 $Y=13332500 $D=9
D1138 gnd! 252 dn PJ=0.0001 m=1 $X=328040 $Y=13542500 $D=9
D1139 252 vdd! dn PJ=0.0002 m=1 $X=330360 $Y=13228100 $D=9
D1140 252 vdd! dn PJ=0.0002 m=1 $X=330360 $Y=13438100 $D=9
D1141 gnd! 252 dn PJ=0.0002 m=1 $X=332680 $Y=13232500 $D=9
D1142 gnd! 252 dn PJ=0.0002 m=1 $X=332680 $Y=13442500 $D=9
D1143 252 vdd! dn PJ=0.0002 m=1 $X=335000 $Y=13228100 $D=9
D1144 252 vdd! dn PJ=0.0002 m=1 $X=335000 $Y=13438100 $D=9
D1145 gnd! A0 dn PJ=0.0002 m=1 $X=1804000 $Y=13232500 $D=9
D1146 gnd! A0 dn PJ=0.0002 m=1 $X=1804000 $Y=13442500 $D=9
D1147 A0 vdd! dn PJ=0.0002 m=1 $X=1806320 $Y=13228100 $D=9
D1148 A0 vdd! dn PJ=0.0002 m=1 $X=1806320 $Y=13438100 $D=9
D1149 gnd! A0 dn PJ=0.0002 m=1 $X=1808640 $Y=13232500 $D=9
D1150 gnd! A0 dn PJ=0.0002 m=1 $X=1808640 $Y=13442500 $D=9
D1151 A0 vdd! dn PJ=0.0001 m=1 $X=1810960 $Y=13228100 $D=9
D1152 A0 vdd! dn PJ=0.0001 m=1 $X=1810960 $Y=13438100 $D=9
D1153 gnd! A0 dn PJ=0.0001 m=1 $X=1814140 $Y=13332500 $D=9
D1154 gnd! A0 dn PJ=0.0001 m=1 $X=1814140 $Y=13542500 $D=9
D1155 A0 vdd! dn PJ=0.0002 m=1 $X=1816460 $Y=13228100 $D=9
D1156 A0 vdd! dn PJ=0.0002 m=1 $X=1816460 $Y=13438100 $D=9
D1157 gnd! A0 dn PJ=0.0002 m=1 $X=1818780 $Y=13232500 $D=9
D1158 gnd! A0 dn PJ=0.0002 m=1 $X=1818780 $Y=13442500 $D=9
D1159 A0 vdd! dn PJ=0.0002 m=1 $X=1821100 $Y=13228100 $D=9
D1160 A0 vdd! dn PJ=0.0002 m=1 $X=1821100 $Y=13438100 $D=9
D1161 gnd! A0 dn PJ=0.0002 m=1 $X=1823420 $Y=13232500 $D=9
D1162 gnd! A0 dn PJ=0.0002 m=1 $X=1823420 $Y=13442500 $D=9
D1163 A0 vdd! dn PJ=0.0001 m=1 $X=1825740 $Y=13228100 $D=9
D1164 A0 vdd! dn PJ=0.0001 m=1 $X=1825740 $Y=13438100 $D=9
D1165 gnd! A0 dn PJ=0.0001 m=1 $X=1828920 $Y=13332500 $D=9
D1166 gnd! A0 dn PJ=0.0001 m=1 $X=1828920 $Y=13542500 $D=9
D1167 A0 vdd! dn PJ=0.0002 m=1 $X=1831240 $Y=13228100 $D=9
D1168 A0 vdd! dn PJ=0.0002 m=1 $X=1831240 $Y=13438100 $D=9
D1169 gnd! A0 dn PJ=0.0002 m=1 $X=1833560 $Y=13232500 $D=9
D1170 gnd! A0 dn PJ=0.0002 m=1 $X=1833560 $Y=13442500 $D=9
D1171 A0 vdd! dn PJ=0.0002 m=1 $X=1835880 $Y=13228100 $D=9
D1172 A0 vdd! dn PJ=0.0002 m=1 $X=1835880 $Y=13438100 $D=9
D1173 gnd! A0 dn PJ=0.0002 m=1 $X=1838200 $Y=13232500 $D=9
D1174 gnd! A0 dn PJ=0.0002 m=1 $X=1838200 $Y=13442500 $D=9
D1175 A0 vdd! dn PJ=0.0001 m=1 $X=1840520 $Y=13228100 $D=9
D1176 A0 vdd! dn PJ=0.0001 m=1 $X=1840520 $Y=13438100 $D=9
D1177 gnd! A0 dn PJ=0.0001 m=1 $X=1843700 $Y=13332500 $D=9
D1178 gnd! A0 dn PJ=0.0001 m=1 $X=1843700 $Y=13542500 $D=9
D1179 A0 vdd! dn PJ=0.0002 m=1 $X=1846020 $Y=13228100 $D=9
D1180 A0 vdd! dn PJ=0.0002 m=1 $X=1846020 $Y=13438100 $D=9
D1181 gnd! A0 dn PJ=0.0002 m=1 $X=1848340 $Y=13232500 $D=9
D1182 gnd! A0 dn PJ=0.0002 m=1 $X=1848340 $Y=13442500 $D=9
D1183 A0 vdd! dn PJ=0.0002 m=1 $X=1850660 $Y=13228100 $D=9
D1184 A0 vdd! dn PJ=0.0002 m=1 $X=1850660 $Y=13438100 $D=9
D1185 gnd! A0 dn PJ=0.0002 m=1 $X=1852980 $Y=13232500 $D=9
D1186 gnd! A0 dn PJ=0.0002 m=1 $X=1852980 $Y=13442500 $D=9
D1187 A0 vdd! dn PJ=0.0001 m=1 $X=1855300 $Y=13228100 $D=9
D1188 A0 vdd! dn PJ=0.0001 m=1 $X=1855300 $Y=13438100 $D=9
D1189 gnd! A0 dn PJ=0.0001 m=1 $X=1858480 $Y=13332500 $D=9
D1190 gnd! A0 dn PJ=0.0001 m=1 $X=1858480 $Y=13542500 $D=9
D1191 A0 vdd! dn PJ=0.0002 m=1 $X=1860800 $Y=13228100 $D=9
D1192 A0 vdd! dn PJ=0.0002 m=1 $X=1860800 $Y=13438100 $D=9
D1193 gnd! A0 dn PJ=0.0002 m=1 $X=1863120 $Y=13232500 $D=9
D1194 gnd! A0 dn PJ=0.0002 m=1 $X=1863120 $Y=13442500 $D=9
D1195 A0 vdd! dn PJ=0.0002 m=1 $X=1865440 $Y=13228100 $D=9
D1196 A0 vdd! dn PJ=0.0002 m=1 $X=1865440 $Y=13438100 $D=9
D1197 gnd! A0 dn PJ=0.0002 m=1 $X=1867760 $Y=13232500 $D=9
D1198 gnd! A0 dn PJ=0.0002 m=1 $X=1867760 $Y=13442500 $D=9
D1199 A0 vdd! dn PJ=0.0001 m=1 $X=1870080 $Y=13228100 $D=9
D1200 A0 vdd! dn PJ=0.0001 m=1 $X=1870080 $Y=13438100 $D=9
D1201 gnd! A0 dn PJ=0.0001 m=1 $X=1873260 $Y=13332500 $D=9
D1202 gnd! A0 dn PJ=0.0001 m=1 $X=1873260 $Y=13542500 $D=9
D1203 A0 vdd! dn PJ=0.0002 m=1 $X=1875580 $Y=13228100 $D=9
D1204 A0 vdd! dn PJ=0.0002 m=1 $X=1875580 $Y=13438100 $D=9
D1205 gnd! A0 dn PJ=0.0002 m=1 $X=1877900 $Y=13232500 $D=9
D1206 gnd! A0 dn PJ=0.0002 m=1 $X=1877900 $Y=13442500 $D=9
D1207 A0 vdd! dn PJ=0.0002 m=1 $X=1880220 $Y=13228100 $D=9
D1208 A0 vdd! dn PJ=0.0002 m=1 $X=1880220 $Y=13438100 $D=9
D1209 gnd! A0 dn PJ=0.0002 m=1 $X=1882540 $Y=13232500 $D=9
D1210 gnd! A0 dn PJ=0.0002 m=1 $X=1882540 $Y=13442500 $D=9
D1211 A0 vdd! dn PJ=0.0001 m=1 $X=1884860 $Y=13228100 $D=9
D1212 A0 vdd! dn PJ=0.0001 m=1 $X=1884860 $Y=13438100 $D=9
D1213 gnd! A0 dn PJ=0.0001 m=1 $X=1888040 $Y=13332500 $D=9
D1214 gnd! A0 dn PJ=0.0001 m=1 $X=1888040 $Y=13542500 $D=9
D1215 A0 vdd! dn PJ=0.0002 m=1 $X=1890360 $Y=13228100 $D=9
D1216 A0 vdd! dn PJ=0.0002 m=1 $X=1890360 $Y=13438100 $D=9
D1217 gnd! A0 dn PJ=0.0002 m=1 $X=1892680 $Y=13232500 $D=9
D1218 gnd! A0 dn PJ=0.0002 m=1 $X=1892680 $Y=13442500 $D=9
D1219 A0 vdd! dn PJ=0.0002 m=1 $X=1895000 $Y=13228100 $D=9
D1220 A0 vdd! dn PJ=0.0002 m=1 $X=1895000 $Y=13438100 $D=9
D1221 gnd! A1 dn PJ=0.0002 m=1 $X=2064000 $Y=13232500 $D=9
D1222 gnd! A1 dn PJ=0.0002 m=1 $X=2064000 $Y=13442500 $D=9
D1223 A1 vdd! dn PJ=0.0002 m=1 $X=2066320 $Y=13228100 $D=9
D1224 A1 vdd! dn PJ=0.0002 m=1 $X=2066320 $Y=13438100 $D=9
D1225 gnd! A1 dn PJ=0.0002 m=1 $X=2068640 $Y=13232500 $D=9
D1226 gnd! A1 dn PJ=0.0002 m=1 $X=2068640 $Y=13442500 $D=9
D1227 A1 vdd! dn PJ=0.0001 m=1 $X=2070960 $Y=13228100 $D=9
D1228 A1 vdd! dn PJ=0.0001 m=1 $X=2070960 $Y=13438100 $D=9
D1229 gnd! A1 dn PJ=0.0001 m=1 $X=2074140 $Y=13332500 $D=9
D1230 gnd! A1 dn PJ=0.0001 m=1 $X=2074140 $Y=13542500 $D=9
D1231 A1 vdd! dn PJ=0.0002 m=1 $X=2076460 $Y=13228100 $D=9
D1232 A1 vdd! dn PJ=0.0002 m=1 $X=2076460 $Y=13438100 $D=9
D1233 gnd! A1 dn PJ=0.0002 m=1 $X=2078780 $Y=13232500 $D=9
D1234 gnd! A1 dn PJ=0.0002 m=1 $X=2078780 $Y=13442500 $D=9
D1235 A1 vdd! dn PJ=0.0002 m=1 $X=2081100 $Y=13228100 $D=9
D1236 A1 vdd! dn PJ=0.0002 m=1 $X=2081100 $Y=13438100 $D=9
D1237 gnd! A1 dn PJ=0.0002 m=1 $X=2083420 $Y=13232500 $D=9
D1238 gnd! A1 dn PJ=0.0002 m=1 $X=2083420 $Y=13442500 $D=9
D1239 A1 vdd! dn PJ=0.0001 m=1 $X=2085740 $Y=13228100 $D=9
D1240 A1 vdd! dn PJ=0.0001 m=1 $X=2085740 $Y=13438100 $D=9
D1241 gnd! A1 dn PJ=0.0001 m=1 $X=2088920 $Y=13332500 $D=9
D1242 gnd! A1 dn PJ=0.0001 m=1 $X=2088920 $Y=13542500 $D=9
D1243 A1 vdd! dn PJ=0.0002 m=1 $X=2091240 $Y=13228100 $D=9
D1244 A1 vdd! dn PJ=0.0002 m=1 $X=2091240 $Y=13438100 $D=9
D1245 gnd! A1 dn PJ=0.0002 m=1 $X=2093560 $Y=13232500 $D=9
D1246 gnd! A1 dn PJ=0.0002 m=1 $X=2093560 $Y=13442500 $D=9
D1247 A1 vdd! dn PJ=0.0002 m=1 $X=2095880 $Y=13228100 $D=9
D1248 A1 vdd! dn PJ=0.0002 m=1 $X=2095880 $Y=13438100 $D=9
D1249 gnd! A1 dn PJ=0.0002 m=1 $X=2098200 $Y=13232500 $D=9
D1250 gnd! A1 dn PJ=0.0002 m=1 $X=2098200 $Y=13442500 $D=9
D1251 A1 vdd! dn PJ=0.0001 m=1 $X=2100520 $Y=13228100 $D=9
D1252 A1 vdd! dn PJ=0.0001 m=1 $X=2100520 $Y=13438100 $D=9
D1253 gnd! A1 dn PJ=0.0001 m=1 $X=2103700 $Y=13332500 $D=9
D1254 gnd! A1 dn PJ=0.0001 m=1 $X=2103700 $Y=13542500 $D=9
D1255 A1 vdd! dn PJ=0.0002 m=1 $X=2106020 $Y=13228100 $D=9
D1256 A1 vdd! dn PJ=0.0002 m=1 $X=2106020 $Y=13438100 $D=9
D1257 gnd! A1 dn PJ=0.0002 m=1 $X=2108340 $Y=13232500 $D=9
D1258 gnd! A1 dn PJ=0.0002 m=1 $X=2108340 $Y=13442500 $D=9
D1259 A1 vdd! dn PJ=0.0002 m=1 $X=2110660 $Y=13228100 $D=9
D1260 A1 vdd! dn PJ=0.0002 m=1 $X=2110660 $Y=13438100 $D=9
D1261 gnd! A1 dn PJ=0.0002 m=1 $X=2112980 $Y=13232500 $D=9
D1262 gnd! A1 dn PJ=0.0002 m=1 $X=2112980 $Y=13442500 $D=9
D1263 A1 vdd! dn PJ=0.0001 m=1 $X=2115300 $Y=13228100 $D=9
D1264 A1 vdd! dn PJ=0.0001 m=1 $X=2115300 $Y=13438100 $D=9
D1265 gnd! A1 dn PJ=0.0001 m=1 $X=2118480 $Y=13332500 $D=9
D1266 gnd! A1 dn PJ=0.0001 m=1 $X=2118480 $Y=13542500 $D=9
D1267 A1 vdd! dn PJ=0.0002 m=1 $X=2120800 $Y=13228100 $D=9
D1268 A1 vdd! dn PJ=0.0002 m=1 $X=2120800 $Y=13438100 $D=9
D1269 gnd! A1 dn PJ=0.0002 m=1 $X=2123120 $Y=13232500 $D=9
D1270 gnd! A1 dn PJ=0.0002 m=1 $X=2123120 $Y=13442500 $D=9
D1271 A1 vdd! dn PJ=0.0002 m=1 $X=2125440 $Y=13228100 $D=9
D1272 A1 vdd! dn PJ=0.0002 m=1 $X=2125440 $Y=13438100 $D=9
D1273 gnd! A1 dn PJ=0.0002 m=1 $X=2127760 $Y=13232500 $D=9
D1274 gnd! A1 dn PJ=0.0002 m=1 $X=2127760 $Y=13442500 $D=9
D1275 A1 vdd! dn PJ=0.0001 m=1 $X=2130080 $Y=13228100 $D=9
D1276 A1 vdd! dn PJ=0.0001 m=1 $X=2130080 $Y=13438100 $D=9
D1277 gnd! A1 dn PJ=0.0001 m=1 $X=2133260 $Y=13332500 $D=9
D1278 gnd! A1 dn PJ=0.0001 m=1 $X=2133260 $Y=13542500 $D=9
D1279 A1 vdd! dn PJ=0.0002 m=1 $X=2135580 $Y=13228100 $D=9
D1280 A1 vdd! dn PJ=0.0002 m=1 $X=2135580 $Y=13438100 $D=9
D1281 gnd! A1 dn PJ=0.0002 m=1 $X=2137900 $Y=13232500 $D=9
D1282 gnd! A1 dn PJ=0.0002 m=1 $X=2137900 $Y=13442500 $D=9
D1283 A1 vdd! dn PJ=0.0002 m=1 $X=2140220 $Y=13228100 $D=9
D1284 A1 vdd! dn PJ=0.0002 m=1 $X=2140220 $Y=13438100 $D=9
D1285 gnd! A1 dn PJ=0.0002 m=1 $X=2142540 $Y=13232500 $D=9
D1286 gnd! A1 dn PJ=0.0002 m=1 $X=2142540 $Y=13442500 $D=9
D1287 A1 vdd! dn PJ=0.0001 m=1 $X=2144860 $Y=13228100 $D=9
D1288 A1 vdd! dn PJ=0.0001 m=1 $X=2144860 $Y=13438100 $D=9
D1289 gnd! A1 dn PJ=0.0001 m=1 $X=2148040 $Y=13332500 $D=9
D1290 gnd! A1 dn PJ=0.0001 m=1 $X=2148040 $Y=13542500 $D=9
D1291 A1 vdd! dn PJ=0.0002 m=1 $X=2150360 $Y=13228100 $D=9
D1292 A1 vdd! dn PJ=0.0002 m=1 $X=2150360 $Y=13438100 $D=9
D1293 gnd! A1 dn PJ=0.0002 m=1 $X=2152680 $Y=13232500 $D=9
D1294 gnd! A1 dn PJ=0.0002 m=1 $X=2152680 $Y=13442500 $D=9
D1295 A1 vdd! dn PJ=0.0002 m=1 $X=2155000 $Y=13228100 $D=9
D1296 A1 vdd! dn PJ=0.0002 m=1 $X=2155000 $Y=13438100 $D=9
D1297 gnd! A3 dn PJ=0.0002 m=1 $X=2584000 $Y=13232500 $D=9
D1298 gnd! A3 dn PJ=0.0002 m=1 $X=2584000 $Y=13442500 $D=9
D1299 A3 vdd! dn PJ=0.0002 m=1 $X=2586320 $Y=13228100 $D=9
D1300 A3 vdd! dn PJ=0.0002 m=1 $X=2586320 $Y=13438100 $D=9
D1301 gnd! A3 dn PJ=0.0002 m=1 $X=2588640 $Y=13232500 $D=9
D1302 gnd! A3 dn PJ=0.0002 m=1 $X=2588640 $Y=13442500 $D=9
D1303 A3 vdd! dn PJ=0.0001 m=1 $X=2590960 $Y=13228100 $D=9
D1304 A3 vdd! dn PJ=0.0001 m=1 $X=2590960 $Y=13438100 $D=9
D1305 gnd! A3 dn PJ=0.0001 m=1 $X=2594140 $Y=13332500 $D=9
D1306 gnd! A3 dn PJ=0.0001 m=1 $X=2594140 $Y=13542500 $D=9
D1307 A3 vdd! dn PJ=0.0002 m=1 $X=2596460 $Y=13228100 $D=9
D1308 A3 vdd! dn PJ=0.0002 m=1 $X=2596460 $Y=13438100 $D=9
D1309 gnd! A3 dn PJ=0.0002 m=1 $X=2598780 $Y=13232500 $D=9
D1310 gnd! A3 dn PJ=0.0002 m=1 $X=2598780 $Y=13442500 $D=9
D1311 A3 vdd! dn PJ=0.0002 m=1 $X=2601100 $Y=13228100 $D=9
D1312 A3 vdd! dn PJ=0.0002 m=1 $X=2601100 $Y=13438100 $D=9
D1313 gnd! A3 dn PJ=0.0002 m=1 $X=2603420 $Y=13232500 $D=9
D1314 gnd! A3 dn PJ=0.0002 m=1 $X=2603420 $Y=13442500 $D=9
D1315 A3 vdd! dn PJ=0.0001 m=1 $X=2605740 $Y=13228100 $D=9
D1316 A3 vdd! dn PJ=0.0001 m=1 $X=2605740 $Y=13438100 $D=9
D1317 gnd! A3 dn PJ=0.0001 m=1 $X=2608920 $Y=13332500 $D=9
D1318 gnd! A3 dn PJ=0.0001 m=1 $X=2608920 $Y=13542500 $D=9
D1319 A3 vdd! dn PJ=0.0002 m=1 $X=2611240 $Y=13228100 $D=9
D1320 A3 vdd! dn PJ=0.0002 m=1 $X=2611240 $Y=13438100 $D=9
D1321 gnd! A3 dn PJ=0.0002 m=1 $X=2613560 $Y=13232500 $D=9
D1322 gnd! A3 dn PJ=0.0002 m=1 $X=2613560 $Y=13442500 $D=9
D1323 A3 vdd! dn PJ=0.0002 m=1 $X=2615880 $Y=13228100 $D=9
D1324 A3 vdd! dn PJ=0.0002 m=1 $X=2615880 $Y=13438100 $D=9
D1325 gnd! A3 dn PJ=0.0002 m=1 $X=2618200 $Y=13232500 $D=9
D1326 gnd! A3 dn PJ=0.0002 m=1 $X=2618200 $Y=13442500 $D=9
D1327 A3 vdd! dn PJ=0.0001 m=1 $X=2620520 $Y=13228100 $D=9
D1328 A3 vdd! dn PJ=0.0001 m=1 $X=2620520 $Y=13438100 $D=9
D1329 gnd! A3 dn PJ=0.0001 m=1 $X=2623700 $Y=13332500 $D=9
D1330 gnd! A3 dn PJ=0.0001 m=1 $X=2623700 $Y=13542500 $D=9
D1331 A3 vdd! dn PJ=0.0002 m=1 $X=2626020 $Y=13228100 $D=9
D1332 A3 vdd! dn PJ=0.0002 m=1 $X=2626020 $Y=13438100 $D=9
D1333 gnd! A3 dn PJ=0.0002 m=1 $X=2628340 $Y=13232500 $D=9
D1334 gnd! A3 dn PJ=0.0002 m=1 $X=2628340 $Y=13442500 $D=9
D1335 A3 vdd! dn PJ=0.0002 m=1 $X=2630660 $Y=13228100 $D=9
D1336 A3 vdd! dn PJ=0.0002 m=1 $X=2630660 $Y=13438100 $D=9
D1337 gnd! A3 dn PJ=0.0002 m=1 $X=2632980 $Y=13232500 $D=9
D1338 gnd! A3 dn PJ=0.0002 m=1 $X=2632980 $Y=13442500 $D=9
D1339 A3 vdd! dn PJ=0.0001 m=1 $X=2635300 $Y=13228100 $D=9
D1340 A3 vdd! dn PJ=0.0001 m=1 $X=2635300 $Y=13438100 $D=9
D1341 gnd! A3 dn PJ=0.0001 m=1 $X=2638480 $Y=13332500 $D=9
D1342 gnd! A3 dn PJ=0.0001 m=1 $X=2638480 $Y=13542500 $D=9
D1343 A3 vdd! dn PJ=0.0002 m=1 $X=2640800 $Y=13228100 $D=9
D1344 A3 vdd! dn PJ=0.0002 m=1 $X=2640800 $Y=13438100 $D=9
D1345 gnd! A3 dn PJ=0.0002 m=1 $X=2643120 $Y=13232500 $D=9
D1346 gnd! A3 dn PJ=0.0002 m=1 $X=2643120 $Y=13442500 $D=9
D1347 A3 vdd! dn PJ=0.0002 m=1 $X=2645440 $Y=13228100 $D=9
D1348 A3 vdd! dn PJ=0.0002 m=1 $X=2645440 $Y=13438100 $D=9
D1349 gnd! A3 dn PJ=0.0002 m=1 $X=2647760 $Y=13232500 $D=9
D1350 gnd! A3 dn PJ=0.0002 m=1 $X=2647760 $Y=13442500 $D=9
D1351 A3 vdd! dn PJ=0.0001 m=1 $X=2650080 $Y=13228100 $D=9
D1352 A3 vdd! dn PJ=0.0001 m=1 $X=2650080 $Y=13438100 $D=9
D1353 gnd! A3 dn PJ=0.0001 m=1 $X=2653260 $Y=13332500 $D=9
D1354 gnd! A3 dn PJ=0.0001 m=1 $X=2653260 $Y=13542500 $D=9
D1355 A3 vdd! dn PJ=0.0002 m=1 $X=2655580 $Y=13228100 $D=9
D1356 A3 vdd! dn PJ=0.0002 m=1 $X=2655580 $Y=13438100 $D=9
D1357 gnd! A3 dn PJ=0.0002 m=1 $X=2657900 $Y=13232500 $D=9
D1358 gnd! A3 dn PJ=0.0002 m=1 $X=2657900 $Y=13442500 $D=9
D1359 A3 vdd! dn PJ=0.0002 m=1 $X=2660220 $Y=13228100 $D=9
D1360 A3 vdd! dn PJ=0.0002 m=1 $X=2660220 $Y=13438100 $D=9
D1361 gnd! A3 dn PJ=0.0002 m=1 $X=2662540 $Y=13232500 $D=9
D1362 gnd! A3 dn PJ=0.0002 m=1 $X=2662540 $Y=13442500 $D=9
D1363 A3 vdd! dn PJ=0.0001 m=1 $X=2664860 $Y=13228100 $D=9
D1364 A3 vdd! dn PJ=0.0001 m=1 $X=2664860 $Y=13438100 $D=9
D1365 gnd! A3 dn PJ=0.0001 m=1 $X=2668040 $Y=13332500 $D=9
D1366 gnd! A3 dn PJ=0.0001 m=1 $X=2668040 $Y=13542500 $D=9
D1367 A3 vdd! dn PJ=0.0002 m=1 $X=2670360 $Y=13228100 $D=9
D1368 A3 vdd! dn PJ=0.0002 m=1 $X=2670360 $Y=13438100 $D=9
D1369 gnd! A3 dn PJ=0.0002 m=1 $X=2672680 $Y=13232500 $D=9
D1370 gnd! A3 dn PJ=0.0002 m=1 $X=2672680 $Y=13442500 $D=9
D1371 A3 vdd! dn PJ=0.0002 m=1 $X=2675000 $Y=13228100 $D=9
D1372 A3 vdd! dn PJ=0.0002 m=1 $X=2675000 $Y=13438100 $D=9
D1373 GND_PAD! VDD_PAD! dn PJ=0.00041 m=1 $X=3254760 $Y=80300 $D=9
D1374 VDD_PAD! vdd! dn PJ=0.00041 m=1 $X=3257260 $Y=80300 $D=9
D1375 vdd! VDD_PAD! dn PJ=0.00041 m=1 $X=3259760 $Y=80300 $D=9
D1376 GND_PAD! VDD_PAD! dn PJ=0.00041 m=1 $X=3264760 $Y=80300 $D=9
D1377 VDD_PAD! vdd! dn PJ=0.00041 m=1 $X=3267260 $Y=80300 $D=9
D1378 vdd! VDD_PAD! dn PJ=0.00041 m=1 $X=3269760 $Y=80300 $D=9
D1379 GND_PAD! VDD_PAD! dn PJ=0.00041 m=1 $X=3274760 $Y=80300 $D=9
D1380 VDD_PAD! vdd! dn PJ=0.00041 m=1 $X=3277260 $Y=80300 $D=9
D1381 vdd! VDD_PAD! dn PJ=0.00041 m=1 $X=3279760 $Y=80300 $D=9
D1382 GND_PAD! VDD_PAD! dn PJ=0.00041 m=1 $X=3284760 $Y=80300 $D=9
D1383 VDD_PAD! vdd! dn PJ=0.00041 m=1 $X=3287260 $Y=80300 $D=9
D1384 vdd! VDD_PAD! dn PJ=0.00041 m=1 $X=3289760 $Y=80300 $D=9
D1385 GND_PAD! VDD_PAD! dn PJ=0.00041 m=1 $X=3294760 $Y=80300 $D=9
D1386 VDD_PAD! vdd! dn PJ=0.00041 m=1 $X=3297260 $Y=80300 $D=9
D1387 vdd! VDD_PAD! dn PJ=0.00041 m=1 $X=3299760 $Y=80300 $D=9
D1388 GND_PAD! VDD_PAD! dn PJ=0.00041 m=1 $X=3304760 $Y=80300 $D=9
D1389 VDD_PAD! vdd! dn PJ=0.00041 m=1 $X=3307260 $Y=80300 $D=9
D1390 vdd! VDD_PAD! dn PJ=0.00041 m=1 $X=3309760 $Y=80300 $D=9
D1391 GND_PAD! VDD_PAD! dn PJ=0.00041 m=1 $X=3314760 $Y=80300 $D=9
D1392 VDD_PAD! vdd! dn PJ=0.00041 m=1 $X=3317260 $Y=80300 $D=9
D1393 vdd! VDD_PAD! dn PJ=0.00041 m=1 $X=3319760 $Y=80300 $D=9
D1394 GND_PAD! VDD_PAD! dn PJ=0.00041 m=1 $X=3324760 $Y=80300 $D=9
D1395 VDD_PAD! vdd! dn PJ=0.00041 m=1 $X=3327260 $Y=80300 $D=9
D1396 vdd! VDD_PAD! dn PJ=0.00041 m=1 $X=3329760 $Y=80300 $D=9
D1397 GND_PAD! VDD_PAD! dn PJ=0.00041 m=1 $X=3334760 $Y=80300 $D=9
D1398 VDD_PAD! vdd! dn PJ=0.00041 m=1 $X=3337260 $Y=80300 $D=9
D1399 vdd! VDD_PAD! dn PJ=0.00041 m=1 $X=3339760 $Y=80300 $D=9
D1400 GND_PAD! VDD_PAD! dn PJ=0.00041 m=1 $X=3344760 $Y=80300 $D=9
D1401 VDD_PAD! vdd! dn PJ=0.00041 m=1 $X=3347260 $Y=80300 $D=9
D1402 gnd! A4 dn PJ=0.0002 m=1 $X=3364000 $Y=13232500 $D=9
D1403 gnd! A4 dn PJ=0.0002 m=1 $X=3364000 $Y=13442500 $D=9
D1404 A4 vdd! dn PJ=0.0002 m=1 $X=3366320 $Y=13228100 $D=9
D1405 A4 vdd! dn PJ=0.0002 m=1 $X=3366320 $Y=13438100 $D=9
D1406 gnd! A4 dn PJ=0.0002 m=1 $X=3368640 $Y=13232500 $D=9
D1407 gnd! A4 dn PJ=0.0002 m=1 $X=3368640 $Y=13442500 $D=9
D1408 A4 vdd! dn PJ=0.0001 m=1 $X=3370960 $Y=13228100 $D=9
D1409 A4 vdd! dn PJ=0.0001 m=1 $X=3370960 $Y=13438100 $D=9
D1410 gnd! A4 dn PJ=0.0001 m=1 $X=3374140 $Y=13332500 $D=9
D1411 gnd! A4 dn PJ=0.0001 m=1 $X=3374140 $Y=13542500 $D=9
D1412 A4 vdd! dn PJ=0.0002 m=1 $X=3376460 $Y=13228100 $D=9
D1413 A4 vdd! dn PJ=0.0002 m=1 $X=3376460 $Y=13438100 $D=9
D1414 gnd! A4 dn PJ=0.0002 m=1 $X=3378780 $Y=13232500 $D=9
D1415 gnd! A4 dn PJ=0.0002 m=1 $X=3378780 $Y=13442500 $D=9
D1416 A4 vdd! dn PJ=0.0002 m=1 $X=3381100 $Y=13228100 $D=9
D1417 A4 vdd! dn PJ=0.0002 m=1 $X=3381100 $Y=13438100 $D=9
D1418 gnd! A4 dn PJ=0.0002 m=1 $X=3383420 $Y=13232500 $D=9
D1419 gnd! A4 dn PJ=0.0002 m=1 $X=3383420 $Y=13442500 $D=9
D1420 A4 vdd! dn PJ=0.0001 m=1 $X=3385740 $Y=13228100 $D=9
D1421 A4 vdd! dn PJ=0.0001 m=1 $X=3385740 $Y=13438100 $D=9
D1422 gnd! A4 dn PJ=0.0001 m=1 $X=3388920 $Y=13332500 $D=9
D1423 gnd! A4 dn PJ=0.0001 m=1 $X=3388920 $Y=13542500 $D=9
D1424 A4 vdd! dn PJ=0.0002 m=1 $X=3391240 $Y=13228100 $D=9
D1425 A4 vdd! dn PJ=0.0002 m=1 $X=3391240 $Y=13438100 $D=9
D1426 gnd! A4 dn PJ=0.0002 m=1 $X=3393560 $Y=13232500 $D=9
D1427 gnd! A4 dn PJ=0.0002 m=1 $X=3393560 $Y=13442500 $D=9
D1428 A4 vdd! dn PJ=0.0002 m=1 $X=3395880 $Y=13228100 $D=9
D1429 A4 vdd! dn PJ=0.0002 m=1 $X=3395880 $Y=13438100 $D=9
D1430 gnd! A4 dn PJ=0.0002 m=1 $X=3398200 $Y=13232500 $D=9
D1431 gnd! A4 dn PJ=0.0002 m=1 $X=3398200 $Y=13442500 $D=9
D1432 A4 vdd! dn PJ=0.0001 m=1 $X=3400520 $Y=13228100 $D=9
D1433 A4 vdd! dn PJ=0.0001 m=1 $X=3400520 $Y=13438100 $D=9
D1434 gnd! A4 dn PJ=0.0001 m=1 $X=3403700 $Y=13332500 $D=9
D1435 gnd! A4 dn PJ=0.0001 m=1 $X=3403700 $Y=13542500 $D=9
D1436 A4 vdd! dn PJ=0.0002 m=1 $X=3406020 $Y=13228100 $D=9
D1437 A4 vdd! dn PJ=0.0002 m=1 $X=3406020 $Y=13438100 $D=9
D1438 gnd! A4 dn PJ=0.0002 m=1 $X=3408340 $Y=13232500 $D=9
D1439 gnd! A4 dn PJ=0.0002 m=1 $X=3408340 $Y=13442500 $D=9
D1440 A4 vdd! dn PJ=0.0002 m=1 $X=3410660 $Y=13228100 $D=9
D1441 A4 vdd! dn PJ=0.0002 m=1 $X=3410660 $Y=13438100 $D=9
D1442 gnd! A4 dn PJ=0.0002 m=1 $X=3412980 $Y=13232500 $D=9
D1443 gnd! A4 dn PJ=0.0002 m=1 $X=3412980 $Y=13442500 $D=9
D1444 A4 vdd! dn PJ=0.0001 m=1 $X=3415300 $Y=13228100 $D=9
D1445 A4 vdd! dn PJ=0.0001 m=1 $X=3415300 $Y=13438100 $D=9
D1446 gnd! A4 dn PJ=0.0001 m=1 $X=3418480 $Y=13332500 $D=9
D1447 gnd! A4 dn PJ=0.0001 m=1 $X=3418480 $Y=13542500 $D=9
D1448 A4 vdd! dn PJ=0.0002 m=1 $X=3420800 $Y=13228100 $D=9
D1449 A4 vdd! dn PJ=0.0002 m=1 $X=3420800 $Y=13438100 $D=9
D1450 gnd! A4 dn PJ=0.0002 m=1 $X=3423120 $Y=13232500 $D=9
D1451 gnd! A4 dn PJ=0.0002 m=1 $X=3423120 $Y=13442500 $D=9
D1452 A4 vdd! dn PJ=0.0002 m=1 $X=3425440 $Y=13228100 $D=9
D1453 A4 vdd! dn PJ=0.0002 m=1 $X=3425440 $Y=13438100 $D=9
D1454 gnd! A4 dn PJ=0.0002 m=1 $X=3427760 $Y=13232500 $D=9
D1455 gnd! A4 dn PJ=0.0002 m=1 $X=3427760 $Y=13442500 $D=9
D1456 A4 vdd! dn PJ=0.0001 m=1 $X=3430080 $Y=13228100 $D=9
D1457 A4 vdd! dn PJ=0.0001 m=1 $X=3430080 $Y=13438100 $D=9
D1458 gnd! A4 dn PJ=0.0001 m=1 $X=3433260 $Y=13332500 $D=9
D1459 gnd! A4 dn PJ=0.0001 m=1 $X=3433260 $Y=13542500 $D=9
D1460 A4 vdd! dn PJ=0.0002 m=1 $X=3435580 $Y=13228100 $D=9
D1461 A4 vdd! dn PJ=0.0002 m=1 $X=3435580 $Y=13438100 $D=9
D1462 gnd! A4 dn PJ=0.0002 m=1 $X=3437900 $Y=13232500 $D=9
D1463 gnd! A4 dn PJ=0.0002 m=1 $X=3437900 $Y=13442500 $D=9
D1464 A4 vdd! dn PJ=0.0002 m=1 $X=3440220 $Y=13228100 $D=9
D1465 A4 vdd! dn PJ=0.0002 m=1 $X=3440220 $Y=13438100 $D=9
D1466 gnd! A4 dn PJ=0.0002 m=1 $X=3442540 $Y=13232500 $D=9
D1467 gnd! A4 dn PJ=0.0002 m=1 $X=3442540 $Y=13442500 $D=9
D1468 A4 vdd! dn PJ=0.0001 m=1 $X=3444860 $Y=13228100 $D=9
D1469 A4 vdd! dn PJ=0.0001 m=1 $X=3444860 $Y=13438100 $D=9
D1470 gnd! A4 dn PJ=0.0001 m=1 $X=3448040 $Y=13332500 $D=9
D1471 gnd! A4 dn PJ=0.0001 m=1 $X=3448040 $Y=13542500 $D=9
D1472 A4 vdd! dn PJ=0.0002 m=1 $X=3450360 $Y=13228100 $D=9
D1473 A4 vdd! dn PJ=0.0002 m=1 $X=3450360 $Y=13438100 $D=9
D1474 gnd! A4 dn PJ=0.0002 m=1 $X=3452680 $Y=13232500 $D=9
D1475 gnd! A4 dn PJ=0.0002 m=1 $X=3452680 $Y=13442500 $D=9
D1476 A4 vdd! dn PJ=0.0002 m=1 $X=3455000 $Y=13228100 $D=9
D1477 A4 vdd! dn PJ=0.0002 m=1 $X=3455000 $Y=13438100 $D=9
D1478 GND_PAD! VDD_PAD! dn PJ=0.00041 m=1 $X=3557480 $Y=80300 $D=9
D1479 GND_PAD! VDD_PAD! dn PJ=0.00041 m=1 $X=3567480 $Y=80300 $D=9
D1480 GND_PAD! VDD_PAD! dn PJ=0.00041 m=1 $X=3577480 $Y=80300 $D=9
D1481 GND_PAD! VDD_PAD! dn PJ=0.00041 m=1 $X=3587480 $Y=80300 $D=9
D1482 GND_PAD! VDD_PAD! dn PJ=0.00041 m=1 $X=3597480 $Y=80300 $D=9
D1483 GND_PAD! VDD_PAD! dn PJ=0.00041 m=1 $X=3607480 $Y=80300 $D=9
D1484 GND_PAD! VDD_PAD! dn PJ=0.00041 m=1 $X=3617480 $Y=80300 $D=9
D1485 GND_PAD! VDD_PAD! dn PJ=0.00041 m=1 $X=3627480 $Y=80300 $D=9
D1486 GND_PAD! VDD_PAD! dn PJ=0.00041 m=1 $X=3637480 $Y=80300 $D=9
D1487 gnd! A6 dn PJ=0.0002 m=1 $X=3884000 $Y=13232500 $D=9
D1488 gnd! A6 dn PJ=0.0002 m=1 $X=3884000 $Y=13442500 $D=9
D1489 A6 vdd! dn PJ=0.0002 m=1 $X=3886320 $Y=13228100 $D=9
D1490 A6 vdd! dn PJ=0.0002 m=1 $X=3886320 $Y=13438100 $D=9
D1491 gnd! A6 dn PJ=0.0002 m=1 $X=3888640 $Y=13232500 $D=9
D1492 gnd! A6 dn PJ=0.0002 m=1 $X=3888640 $Y=13442500 $D=9
D1493 A6 vdd! dn PJ=0.0001 m=1 $X=3890960 $Y=13228100 $D=9
D1494 A6 vdd! dn PJ=0.0001 m=1 $X=3890960 $Y=13438100 $D=9
D1495 gnd! A6 dn PJ=0.0001 m=1 $X=3894140 $Y=13332500 $D=9
D1496 gnd! A6 dn PJ=0.0001 m=1 $X=3894140 $Y=13542500 $D=9
D1497 A6 vdd! dn PJ=0.0002 m=1 $X=3896460 $Y=13228100 $D=9
D1498 A6 vdd! dn PJ=0.0002 m=1 $X=3896460 $Y=13438100 $D=9
D1499 gnd! A6 dn PJ=0.0002 m=1 $X=3898780 $Y=13232500 $D=9
D1500 gnd! A6 dn PJ=0.0002 m=1 $X=3898780 $Y=13442500 $D=9
D1501 A6 vdd! dn PJ=0.0002 m=1 $X=3901100 $Y=13228100 $D=9
D1502 A6 vdd! dn PJ=0.0002 m=1 $X=3901100 $Y=13438100 $D=9
D1503 gnd! A6 dn PJ=0.0002 m=1 $X=3903420 $Y=13232500 $D=9
D1504 gnd! A6 dn PJ=0.0002 m=1 $X=3903420 $Y=13442500 $D=9
D1505 A6 vdd! dn PJ=0.0001 m=1 $X=3905740 $Y=13228100 $D=9
D1506 A6 vdd! dn PJ=0.0001 m=1 $X=3905740 $Y=13438100 $D=9
D1507 gnd! A6 dn PJ=0.0001 m=1 $X=3908920 $Y=13332500 $D=9
D1508 gnd! A6 dn PJ=0.0001 m=1 $X=3908920 $Y=13542500 $D=9
D1509 A6 vdd! dn PJ=0.0002 m=1 $X=3911240 $Y=13228100 $D=9
D1510 A6 vdd! dn PJ=0.0002 m=1 $X=3911240 $Y=13438100 $D=9
D1511 gnd! A6 dn PJ=0.0002 m=1 $X=3913560 $Y=13232500 $D=9
D1512 gnd! A6 dn PJ=0.0002 m=1 $X=3913560 $Y=13442500 $D=9
D1513 A6 vdd! dn PJ=0.0002 m=1 $X=3915880 $Y=13228100 $D=9
D1514 A6 vdd! dn PJ=0.0002 m=1 $X=3915880 $Y=13438100 $D=9
D1515 gnd! A6 dn PJ=0.0002 m=1 $X=3918200 $Y=13232500 $D=9
D1516 gnd! A6 dn PJ=0.0002 m=1 $X=3918200 $Y=13442500 $D=9
D1517 A6 vdd! dn PJ=0.0001 m=1 $X=3920520 $Y=13228100 $D=9
D1518 A6 vdd! dn PJ=0.0001 m=1 $X=3920520 $Y=13438100 $D=9
D1519 gnd! A6 dn PJ=0.0001 m=1 $X=3923700 $Y=13332500 $D=9
D1520 gnd! A6 dn PJ=0.0001 m=1 $X=3923700 $Y=13542500 $D=9
D1521 A6 vdd! dn PJ=0.0002 m=1 $X=3926020 $Y=13228100 $D=9
D1522 A6 vdd! dn PJ=0.0002 m=1 $X=3926020 $Y=13438100 $D=9
D1523 gnd! A6 dn PJ=0.0002 m=1 $X=3928340 $Y=13232500 $D=9
D1524 gnd! A6 dn PJ=0.0002 m=1 $X=3928340 $Y=13442500 $D=9
D1525 A6 vdd! dn PJ=0.0002 m=1 $X=3930660 $Y=13228100 $D=9
D1526 A6 vdd! dn PJ=0.0002 m=1 $X=3930660 $Y=13438100 $D=9
D1527 gnd! A6 dn PJ=0.0002 m=1 $X=3932980 $Y=13232500 $D=9
D1528 gnd! A6 dn PJ=0.0002 m=1 $X=3932980 $Y=13442500 $D=9
D1529 A6 vdd! dn PJ=0.0001 m=1 $X=3935300 $Y=13228100 $D=9
D1530 A6 vdd! dn PJ=0.0001 m=1 $X=3935300 $Y=13438100 $D=9
D1531 gnd! A6 dn PJ=0.0001 m=1 $X=3938480 $Y=13332500 $D=9
D1532 gnd! A6 dn PJ=0.0001 m=1 $X=3938480 $Y=13542500 $D=9
D1533 A6 vdd! dn PJ=0.0002 m=1 $X=3940800 $Y=13228100 $D=9
D1534 A6 vdd! dn PJ=0.0002 m=1 $X=3940800 $Y=13438100 $D=9
D1535 gnd! A6 dn PJ=0.0002 m=1 $X=3943120 $Y=13232500 $D=9
D1536 gnd! A6 dn PJ=0.0002 m=1 $X=3943120 $Y=13442500 $D=9
D1537 A6 vdd! dn PJ=0.0002 m=1 $X=3945440 $Y=13228100 $D=9
D1538 A6 vdd! dn PJ=0.0002 m=1 $X=3945440 $Y=13438100 $D=9
D1539 gnd! A6 dn PJ=0.0002 m=1 $X=3947760 $Y=13232500 $D=9
D1540 gnd! A6 dn PJ=0.0002 m=1 $X=3947760 $Y=13442500 $D=9
D1541 A6 vdd! dn PJ=0.0001 m=1 $X=3950080 $Y=13228100 $D=9
D1542 A6 vdd! dn PJ=0.0001 m=1 $X=3950080 $Y=13438100 $D=9
D1543 gnd! A6 dn PJ=0.0001 m=1 $X=3953260 $Y=13332500 $D=9
D1544 gnd! A6 dn PJ=0.0001 m=1 $X=3953260 $Y=13542500 $D=9
D1545 A6 vdd! dn PJ=0.0002 m=1 $X=3955580 $Y=13228100 $D=9
D1546 A6 vdd! dn PJ=0.0002 m=1 $X=3955580 $Y=13438100 $D=9
D1547 gnd! A6 dn PJ=0.0002 m=1 $X=3957900 $Y=13232500 $D=9
D1548 gnd! A6 dn PJ=0.0002 m=1 $X=3957900 $Y=13442500 $D=9
D1549 A6 vdd! dn PJ=0.0002 m=1 $X=3960220 $Y=13228100 $D=9
D1550 A6 vdd! dn PJ=0.0002 m=1 $X=3960220 $Y=13438100 $D=9
D1551 gnd! A6 dn PJ=0.0002 m=1 $X=3962540 $Y=13232500 $D=9
D1552 gnd! A6 dn PJ=0.0002 m=1 $X=3962540 $Y=13442500 $D=9
D1553 A6 vdd! dn PJ=0.0001 m=1 $X=3964860 $Y=13228100 $D=9
D1554 A6 vdd! dn PJ=0.0001 m=1 $X=3964860 $Y=13438100 $D=9
D1555 gnd! A6 dn PJ=0.0001 m=1 $X=3968040 $Y=13332500 $D=9
D1556 gnd! A6 dn PJ=0.0001 m=1 $X=3968040 $Y=13542500 $D=9
D1557 A6 vdd! dn PJ=0.0002 m=1 $X=3970360 $Y=13228100 $D=9
D1558 A6 vdd! dn PJ=0.0002 m=1 $X=3970360 $Y=13438100 $D=9
D1559 gnd! A6 dn PJ=0.0002 m=1 $X=3972680 $Y=13232500 $D=9
D1560 gnd! A6 dn PJ=0.0002 m=1 $X=3972680 $Y=13442500 $D=9
D1561 A6 vdd! dn PJ=0.0002 m=1 $X=3975000 $Y=13228100 $D=9
D1562 A6 vdd! dn PJ=0.0002 m=1 $X=3975000 $Y=13438100 $D=9
D1563 gnd! A7 dn PJ=0.0002 m=1 $X=4144000 $Y=13232500 $D=9
D1564 gnd! A7 dn PJ=0.0002 m=1 $X=4144000 $Y=13442500 $D=9
D1565 A7 vdd! dn PJ=0.0002 m=1 $X=4146320 $Y=13228100 $D=9
D1566 A7 vdd! dn PJ=0.0002 m=1 $X=4146320 $Y=13438100 $D=9
D1567 gnd! A7 dn PJ=0.0002 m=1 $X=4148640 $Y=13232500 $D=9
D1568 gnd! A7 dn PJ=0.0002 m=1 $X=4148640 $Y=13442500 $D=9
D1569 A7 vdd! dn PJ=0.0001 m=1 $X=4150960 $Y=13228100 $D=9
D1570 A7 vdd! dn PJ=0.0001 m=1 $X=4150960 $Y=13438100 $D=9
D1571 gnd! A7 dn PJ=0.0001 m=1 $X=4154140 $Y=13332500 $D=9
D1572 gnd! A7 dn PJ=0.0001 m=1 $X=4154140 $Y=13542500 $D=9
D1573 A7 vdd! dn PJ=0.0002 m=1 $X=4156460 $Y=13228100 $D=9
D1574 A7 vdd! dn PJ=0.0002 m=1 $X=4156460 $Y=13438100 $D=9
D1575 gnd! A7 dn PJ=0.0002 m=1 $X=4158780 $Y=13232500 $D=9
D1576 gnd! A7 dn PJ=0.0002 m=1 $X=4158780 $Y=13442500 $D=9
D1577 A7 vdd! dn PJ=0.0002 m=1 $X=4161100 $Y=13228100 $D=9
D1578 A7 vdd! dn PJ=0.0002 m=1 $X=4161100 $Y=13438100 $D=9
D1579 gnd! A7 dn PJ=0.0002 m=1 $X=4163420 $Y=13232500 $D=9
D1580 gnd! A7 dn PJ=0.0002 m=1 $X=4163420 $Y=13442500 $D=9
D1581 A7 vdd! dn PJ=0.0001 m=1 $X=4165740 $Y=13228100 $D=9
D1582 A7 vdd! dn PJ=0.0001 m=1 $X=4165740 $Y=13438100 $D=9
D1583 gnd! A7 dn PJ=0.0001 m=1 $X=4168920 $Y=13332500 $D=9
D1584 gnd! A7 dn PJ=0.0001 m=1 $X=4168920 $Y=13542500 $D=9
D1585 A7 vdd! dn PJ=0.0002 m=1 $X=4171240 $Y=13228100 $D=9
D1586 A7 vdd! dn PJ=0.0002 m=1 $X=4171240 $Y=13438100 $D=9
D1587 gnd! A7 dn PJ=0.0002 m=1 $X=4173560 $Y=13232500 $D=9
D1588 gnd! A7 dn PJ=0.0002 m=1 $X=4173560 $Y=13442500 $D=9
D1589 A7 vdd! dn PJ=0.0002 m=1 $X=4175880 $Y=13228100 $D=9
D1590 A7 vdd! dn PJ=0.0002 m=1 $X=4175880 $Y=13438100 $D=9
D1591 gnd! A7 dn PJ=0.0002 m=1 $X=4178200 $Y=13232500 $D=9
D1592 gnd! A7 dn PJ=0.0002 m=1 $X=4178200 $Y=13442500 $D=9
D1593 A7 vdd! dn PJ=0.0001 m=1 $X=4180520 $Y=13228100 $D=9
D1594 A7 vdd! dn PJ=0.0001 m=1 $X=4180520 $Y=13438100 $D=9
D1595 gnd! A7 dn PJ=0.0001 m=1 $X=4183700 $Y=13332500 $D=9
D1596 gnd! A7 dn PJ=0.0001 m=1 $X=4183700 $Y=13542500 $D=9
D1597 A7 vdd! dn PJ=0.0002 m=1 $X=4186020 $Y=13228100 $D=9
D1598 A7 vdd! dn PJ=0.0002 m=1 $X=4186020 $Y=13438100 $D=9
D1599 gnd! A7 dn PJ=0.0002 m=1 $X=4188340 $Y=13232500 $D=9
D1600 gnd! A7 dn PJ=0.0002 m=1 $X=4188340 $Y=13442500 $D=9
D1601 A7 vdd! dn PJ=0.0002 m=1 $X=4190660 $Y=13228100 $D=9
D1602 A7 vdd! dn PJ=0.0002 m=1 $X=4190660 $Y=13438100 $D=9
D1603 gnd! A7 dn PJ=0.0002 m=1 $X=4192980 $Y=13232500 $D=9
D1604 gnd! A7 dn PJ=0.0002 m=1 $X=4192980 $Y=13442500 $D=9
D1605 A7 vdd! dn PJ=0.0001 m=1 $X=4195300 $Y=13228100 $D=9
D1606 A7 vdd! dn PJ=0.0001 m=1 $X=4195300 $Y=13438100 $D=9
D1607 gnd! A7 dn PJ=0.0001 m=1 $X=4198480 $Y=13332500 $D=9
D1608 gnd! A7 dn PJ=0.0001 m=1 $X=4198480 $Y=13542500 $D=9
D1609 A7 vdd! dn PJ=0.0002 m=1 $X=4200800 $Y=13228100 $D=9
D1610 A7 vdd! dn PJ=0.0002 m=1 $X=4200800 $Y=13438100 $D=9
D1611 gnd! A7 dn PJ=0.0002 m=1 $X=4203120 $Y=13232500 $D=9
D1612 gnd! A7 dn PJ=0.0002 m=1 $X=4203120 $Y=13442500 $D=9
D1613 A7 vdd! dn PJ=0.0002 m=1 $X=4205440 $Y=13228100 $D=9
D1614 A7 vdd! dn PJ=0.0002 m=1 $X=4205440 $Y=13438100 $D=9
D1615 gnd! A7 dn PJ=0.0002 m=1 $X=4207760 $Y=13232500 $D=9
D1616 gnd! A7 dn PJ=0.0002 m=1 $X=4207760 $Y=13442500 $D=9
D1617 A7 vdd! dn PJ=0.0001 m=1 $X=4210080 $Y=13228100 $D=9
D1618 A7 vdd! dn PJ=0.0001 m=1 $X=4210080 $Y=13438100 $D=9
D1619 gnd! A7 dn PJ=0.0001 m=1 $X=4213260 $Y=13332500 $D=9
D1620 gnd! A7 dn PJ=0.0001 m=1 $X=4213260 $Y=13542500 $D=9
D1621 A7 vdd! dn PJ=0.0002 m=1 $X=4215580 $Y=13228100 $D=9
D1622 A7 vdd! dn PJ=0.0002 m=1 $X=4215580 $Y=13438100 $D=9
D1623 gnd! A7 dn PJ=0.0002 m=1 $X=4217900 $Y=13232500 $D=9
D1624 gnd! A7 dn PJ=0.0002 m=1 $X=4217900 $Y=13442500 $D=9
D1625 A7 vdd! dn PJ=0.0002 m=1 $X=4220220 $Y=13228100 $D=9
D1626 A7 vdd! dn PJ=0.0002 m=1 $X=4220220 $Y=13438100 $D=9
D1627 gnd! A7 dn PJ=0.0002 m=1 $X=4222540 $Y=13232500 $D=9
D1628 gnd! A7 dn PJ=0.0002 m=1 $X=4222540 $Y=13442500 $D=9
D1629 A7 vdd! dn PJ=0.0001 m=1 $X=4224860 $Y=13228100 $D=9
D1630 A7 vdd! dn PJ=0.0001 m=1 $X=4224860 $Y=13438100 $D=9
D1631 gnd! A7 dn PJ=0.0001 m=1 $X=4228040 $Y=13332500 $D=9
D1632 gnd! A7 dn PJ=0.0001 m=1 $X=4228040 $Y=13542500 $D=9
D1633 A7 vdd! dn PJ=0.0002 m=1 $X=4230360 $Y=13228100 $D=9
D1634 A7 vdd! dn PJ=0.0002 m=1 $X=4230360 $Y=13438100 $D=9
D1635 gnd! A7 dn PJ=0.0002 m=1 $X=4232680 $Y=13232500 $D=9
D1636 gnd! A7 dn PJ=0.0002 m=1 $X=4232680 $Y=13442500 $D=9
D1637 A7 vdd! dn PJ=0.0002 m=1 $X=4235000 $Y=13228100 $D=9
D1638 A7 vdd! dn PJ=0.0002 m=1 $X=4235000 $Y=13438100 $D=9
D1639 gnd! A20 dn PJ=0.0002 m=1 $X=6224000 $Y=13232500 $D=9
D1640 gnd! A20 dn PJ=0.0002 m=1 $X=6224000 $Y=13442500 $D=9
D1641 A20 vdd! dn PJ=0.0002 m=1 $X=6226320 $Y=13228100 $D=9
D1642 A20 vdd! dn PJ=0.0002 m=1 $X=6226320 $Y=13438100 $D=9
D1643 gnd! A20 dn PJ=0.0002 m=1 $X=6228640 $Y=13232500 $D=9
D1644 gnd! A20 dn PJ=0.0002 m=1 $X=6228640 $Y=13442500 $D=9
D1645 A20 vdd! dn PJ=0.0001 m=1 $X=6230960 $Y=13228100 $D=9
D1646 A20 vdd! dn PJ=0.0001 m=1 $X=6230960 $Y=13438100 $D=9
D1647 gnd! A20 dn PJ=0.0001 m=1 $X=6234140 $Y=13332500 $D=9
D1648 gnd! A20 dn PJ=0.0001 m=1 $X=6234140 $Y=13542500 $D=9
D1649 A20 vdd! dn PJ=0.0002 m=1 $X=6236460 $Y=13228100 $D=9
D1650 A20 vdd! dn PJ=0.0002 m=1 $X=6236460 $Y=13438100 $D=9
D1651 gnd! A20 dn PJ=0.0002 m=1 $X=6238780 $Y=13232500 $D=9
D1652 gnd! A20 dn PJ=0.0002 m=1 $X=6238780 $Y=13442500 $D=9
D1653 A20 vdd! dn PJ=0.0002 m=1 $X=6241100 $Y=13228100 $D=9
D1654 A20 vdd! dn PJ=0.0002 m=1 $X=6241100 $Y=13438100 $D=9
D1655 gnd! A20 dn PJ=0.0002 m=1 $X=6243420 $Y=13232500 $D=9
D1656 gnd! A20 dn PJ=0.0002 m=1 $X=6243420 $Y=13442500 $D=9
D1657 A20 vdd! dn PJ=0.0001 m=1 $X=6245740 $Y=13228100 $D=9
D1658 A20 vdd! dn PJ=0.0001 m=1 $X=6245740 $Y=13438100 $D=9
D1659 gnd! A20 dn PJ=0.0001 m=1 $X=6248920 $Y=13332500 $D=9
D1660 gnd! A20 dn PJ=0.0001 m=1 $X=6248920 $Y=13542500 $D=9
D1661 A20 vdd! dn PJ=0.0002 m=1 $X=6251240 $Y=13228100 $D=9
D1662 A20 vdd! dn PJ=0.0002 m=1 $X=6251240 $Y=13438100 $D=9
D1663 gnd! A20 dn PJ=0.0002 m=1 $X=6253560 $Y=13232500 $D=9
D1664 gnd! A20 dn PJ=0.0002 m=1 $X=6253560 $Y=13442500 $D=9
D1665 A20 vdd! dn PJ=0.0002 m=1 $X=6255880 $Y=13228100 $D=9
D1666 A20 vdd! dn PJ=0.0002 m=1 $X=6255880 $Y=13438100 $D=9
D1667 gnd! A20 dn PJ=0.0002 m=1 $X=6258200 $Y=13232500 $D=9
D1668 gnd! A20 dn PJ=0.0002 m=1 $X=6258200 $Y=13442500 $D=9
D1669 A20 vdd! dn PJ=0.0001 m=1 $X=6260520 $Y=13228100 $D=9
D1670 A20 vdd! dn PJ=0.0001 m=1 $X=6260520 $Y=13438100 $D=9
D1671 gnd! A20 dn PJ=0.0001 m=1 $X=6263700 $Y=13332500 $D=9
D1672 gnd! A20 dn PJ=0.0001 m=1 $X=6263700 $Y=13542500 $D=9
D1673 A20 vdd! dn PJ=0.0002 m=1 $X=6266020 $Y=13228100 $D=9
D1674 A20 vdd! dn PJ=0.0002 m=1 $X=6266020 $Y=13438100 $D=9
D1675 gnd! A20 dn PJ=0.0002 m=1 $X=6268340 $Y=13232500 $D=9
D1676 gnd! A20 dn PJ=0.0002 m=1 $X=6268340 $Y=13442500 $D=9
D1677 A20 vdd! dn PJ=0.0002 m=1 $X=6270660 $Y=13228100 $D=9
D1678 A20 vdd! dn PJ=0.0002 m=1 $X=6270660 $Y=13438100 $D=9
D1679 gnd! A20 dn PJ=0.0002 m=1 $X=6272980 $Y=13232500 $D=9
D1680 gnd! A20 dn PJ=0.0002 m=1 $X=6272980 $Y=13442500 $D=9
D1681 A20 vdd! dn PJ=0.0001 m=1 $X=6275300 $Y=13228100 $D=9
D1682 A20 vdd! dn PJ=0.0001 m=1 $X=6275300 $Y=13438100 $D=9
D1683 gnd! A20 dn PJ=0.0001 m=1 $X=6278480 $Y=13332500 $D=9
D1684 gnd! A20 dn PJ=0.0001 m=1 $X=6278480 $Y=13542500 $D=9
D1685 A20 vdd! dn PJ=0.0002 m=1 $X=6280800 $Y=13228100 $D=9
D1686 A20 vdd! dn PJ=0.0002 m=1 $X=6280800 $Y=13438100 $D=9
D1687 gnd! A20 dn PJ=0.0002 m=1 $X=6283120 $Y=13232500 $D=9
D1688 gnd! A20 dn PJ=0.0002 m=1 $X=6283120 $Y=13442500 $D=9
D1689 A20 vdd! dn PJ=0.0002 m=1 $X=6285440 $Y=13228100 $D=9
D1690 A20 vdd! dn PJ=0.0002 m=1 $X=6285440 $Y=13438100 $D=9
D1691 gnd! A20 dn PJ=0.0002 m=1 $X=6287760 $Y=13232500 $D=9
D1692 gnd! A20 dn PJ=0.0002 m=1 $X=6287760 $Y=13442500 $D=9
D1693 A20 vdd! dn PJ=0.0001 m=1 $X=6290080 $Y=13228100 $D=9
D1694 A20 vdd! dn PJ=0.0001 m=1 $X=6290080 $Y=13438100 $D=9
D1695 gnd! A20 dn PJ=0.0001 m=1 $X=6293260 $Y=13332500 $D=9
D1696 gnd! A20 dn PJ=0.0001 m=1 $X=6293260 $Y=13542500 $D=9
D1697 A20 vdd! dn PJ=0.0002 m=1 $X=6295580 $Y=13228100 $D=9
D1698 A20 vdd! dn PJ=0.0002 m=1 $X=6295580 $Y=13438100 $D=9
D1699 gnd! A20 dn PJ=0.0002 m=1 $X=6297900 $Y=13232500 $D=9
D1700 gnd! A20 dn PJ=0.0002 m=1 $X=6297900 $Y=13442500 $D=9
D1701 A20 vdd! dn PJ=0.0002 m=1 $X=6300220 $Y=13228100 $D=9
D1702 A20 vdd! dn PJ=0.0002 m=1 $X=6300220 $Y=13438100 $D=9
D1703 gnd! A20 dn PJ=0.0002 m=1 $X=6302540 $Y=13232500 $D=9
D1704 gnd! A20 dn PJ=0.0002 m=1 $X=6302540 $Y=13442500 $D=9
D1705 A20 vdd! dn PJ=0.0001 m=1 $X=6304860 $Y=13228100 $D=9
D1706 A20 vdd! dn PJ=0.0001 m=1 $X=6304860 $Y=13438100 $D=9
D1707 gnd! A20 dn PJ=0.0001 m=1 $X=6308040 $Y=13332500 $D=9
D1708 gnd! A20 dn PJ=0.0001 m=1 $X=6308040 $Y=13542500 $D=9
D1709 A20 vdd! dn PJ=0.0002 m=1 $X=6310360 $Y=13228100 $D=9
D1710 A20 vdd! dn PJ=0.0002 m=1 $X=6310360 $Y=13438100 $D=9
D1711 gnd! A20 dn PJ=0.0002 m=1 $X=6312680 $Y=13232500 $D=9
D1712 gnd! A20 dn PJ=0.0002 m=1 $X=6312680 $Y=13442500 $D=9
D1713 A20 vdd! dn PJ=0.0002 m=1 $X=6315000 $Y=13228100 $D=9
D1714 A20 vdd! dn PJ=0.0002 m=1 $X=6315000 $Y=13438100 $D=9
D1715 gnd! vdd! dn PJ=0.00041 m=1 $X=7154740 $Y=80300 $D=9
D1716 vdd! VDD_PAD! dn PJ=0.00041 m=1 $X=7157240 $Y=80300 $D=9
D1717 gnd! vdd! dn PJ=0.00041 m=1 $X=7164740 $Y=80300 $D=9
D1718 vdd! VDD_PAD! dn PJ=0.00041 m=1 $X=7167240 $Y=80300 $D=9
D1719 gnd! vdd! dn PJ=0.00041 m=1 $X=7174740 $Y=80300 $D=9
D1720 vdd! VDD_PAD! dn PJ=0.00041 m=1 $X=7177240 $Y=80300 $D=9
D1721 gnd! vdd! dn PJ=0.00041 m=1 $X=7184740 $Y=80300 $D=9
D1722 vdd! VDD_PAD! dn PJ=0.00041 m=1 $X=7187240 $Y=80300 $D=9
D1723 gnd! vdd! dn PJ=0.00041 m=1 $X=7194740 $Y=80300 $D=9
D1724 vdd! VDD_PAD! dn PJ=0.00041 m=1 $X=7197240 $Y=80300 $D=9
D1725 gnd! vdd! dn PJ=0.00041 m=1 $X=7204740 $Y=80300 $D=9
D1726 vdd! VDD_PAD! dn PJ=0.00041 m=1 $X=7207240 $Y=80300 $D=9
D1727 gnd! vdd! dn PJ=0.00041 m=1 $X=7214740 $Y=80300 $D=9
D1728 vdd! VDD_PAD! dn PJ=0.00041 m=1 $X=7217240 $Y=80300 $D=9
D1729 gnd! vdd! dn PJ=0.00041 m=1 $X=7224740 $Y=80300 $D=9
D1730 vdd! VDD_PAD! dn PJ=0.00041 m=1 $X=7227240 $Y=80300 $D=9
D1731 gnd! vdd! dn PJ=0.00041 m=1 $X=7234740 $Y=80300 $D=9
D1732 vdd! VDD_PAD! dn PJ=0.00041 m=1 $X=7237240 $Y=80300 $D=9
D1733 gnd! vdd! dn PJ=0.00041 m=1 $X=7244740 $Y=80300 $D=9
D1734 gnd! vdd! dn PJ=0.00041 m=1 $X=7457460 $Y=80300 $D=9
D1735 vdd! VDD_PAD! dn PJ=0.00041 m=1 $X=7459960 $Y=80300 $D=9
D1736 gnd! vdd! dn PJ=0.00041 m=1 $X=7467460 $Y=80300 $D=9
D1737 vdd! VDD_PAD! dn PJ=0.00041 m=1 $X=7469960 $Y=80300 $D=9
D1738 gnd! vdd! dn PJ=0.00041 m=1 $X=7477460 $Y=80300 $D=9
D1739 vdd! VDD_PAD! dn PJ=0.00041 m=1 $X=7479960 $Y=80300 $D=9
D1740 gnd! vdd! dn PJ=0.00041 m=1 $X=7487460 $Y=80300 $D=9
D1741 vdd! VDD_PAD! dn PJ=0.00041 m=1 $X=7489960 $Y=80300 $D=9
D1742 gnd! vdd! dn PJ=0.00041 m=1 $X=7497460 $Y=80300 $D=9
D1743 vdd! VDD_PAD! dn PJ=0.00041 m=1 $X=7499960 $Y=80300 $D=9
D1744 gnd! vdd! dn PJ=0.00041 m=1 $X=7507460 $Y=80300 $D=9
D1745 vdd! VDD_PAD! dn PJ=0.00041 m=1 $X=7509960 $Y=80300 $D=9
D1746 gnd! vdd! dn PJ=0.00041 m=1 $X=7517460 $Y=80300 $D=9
D1747 vdd! VDD_PAD! dn PJ=0.00041 m=1 $X=7519960 $Y=80300 $D=9
D1748 gnd! vdd! dn PJ=0.00041 m=1 $X=7527460 $Y=80300 $D=9
D1749 vdd! VDD_PAD! dn PJ=0.00041 m=1 $X=7529960 $Y=80300 $D=9
D1750 gnd! vdd! dn PJ=0.00041 m=1 $X=7537460 $Y=80300 $D=9
D1751 vdd! VDD_PAD! dn PJ=0.00041 m=1 $X=7539960 $Y=80300 $D=9
D1752 GND_PAD! VDD_PAD! dn PJ=0.00041 m=1 $X=7754760 $Y=80300 $D=9
D1753 VDD_PAD! vdd! dn PJ=0.00041 m=1 $X=7757260 $Y=80300 $D=9
D1754 vdd! VDD_PAD! dn PJ=0.00041 m=1 $X=7759760 $Y=80300 $D=9
D1755 GND_PAD! VDD_PAD! dn PJ=0.00041 m=1 $X=7764760 $Y=80300 $D=9
D1756 VDD_PAD! vdd! dn PJ=0.00041 m=1 $X=7767260 $Y=80300 $D=9
D1757 vdd! VDD_PAD! dn PJ=0.00041 m=1 $X=7769760 $Y=80300 $D=9
D1758 GND_PAD! VDD_PAD! dn PJ=0.00041 m=1 $X=7774760 $Y=80300 $D=9
D1759 VDD_PAD! vdd! dn PJ=0.00041 m=1 $X=7777260 $Y=80300 $D=9
D1760 vdd! VDD_PAD! dn PJ=0.00041 m=1 $X=7779760 $Y=80300 $D=9
D1761 gnd! CS2 dn PJ=0.0002 m=1 $X=7784000 $Y=13232500 $D=9
D1762 gnd! CS2 dn PJ=0.0002 m=1 $X=7784000 $Y=13442500 $D=9
D1763 GND_PAD! VDD_PAD! dn PJ=0.00041 m=1 $X=7784760 $Y=80300 $D=9
D1764 CS2 vdd! dn PJ=0.0002 m=1 $X=7786320 $Y=13228100 $D=9
D1765 CS2 vdd! dn PJ=0.0002 m=1 $X=7786320 $Y=13438100 $D=9
D1766 VDD_PAD! vdd! dn PJ=0.00041 m=1 $X=7787260 $Y=80300 $D=9
D1767 gnd! CS2 dn PJ=0.0002 m=1 $X=7788640 $Y=13232500 $D=9
D1768 gnd! CS2 dn PJ=0.0002 m=1 $X=7788640 $Y=13442500 $D=9
D1769 vdd! VDD_PAD! dn PJ=0.00041 m=1 $X=7789760 $Y=80300 $D=9
D1770 CS2 vdd! dn PJ=0.0001 m=1 $X=7790960 $Y=13228100 $D=9
D1771 CS2 vdd! dn PJ=0.0001 m=1 $X=7790960 $Y=13438100 $D=9
D1772 gnd! CS2 dn PJ=0.0001 m=1 $X=7794140 $Y=13332500 $D=9
D1773 gnd! CS2 dn PJ=0.0001 m=1 $X=7794140 $Y=13542500 $D=9
D1774 GND_PAD! VDD_PAD! dn PJ=0.00041 m=1 $X=7794760 $Y=80300 $D=9
D1775 CS2 vdd! dn PJ=0.0002 m=1 $X=7796460 $Y=13228100 $D=9
D1776 CS2 vdd! dn PJ=0.0002 m=1 $X=7796460 $Y=13438100 $D=9
D1777 VDD_PAD! vdd! dn PJ=0.00041 m=1 $X=7797260 $Y=80300 $D=9
D1778 gnd! CS2 dn PJ=0.0002 m=1 $X=7798780 $Y=13232500 $D=9
D1779 gnd! CS2 dn PJ=0.0002 m=1 $X=7798780 $Y=13442500 $D=9
D1780 vdd! VDD_PAD! dn PJ=0.00041 m=1 $X=7799760 $Y=80300 $D=9
D1781 CS2 vdd! dn PJ=0.0002 m=1 $X=7801100 $Y=13228100 $D=9
D1782 CS2 vdd! dn PJ=0.0002 m=1 $X=7801100 $Y=13438100 $D=9
D1783 gnd! CS2 dn PJ=0.0002 m=1 $X=7803420 $Y=13232500 $D=9
D1784 gnd! CS2 dn PJ=0.0002 m=1 $X=7803420 $Y=13442500 $D=9
D1785 GND_PAD! VDD_PAD! dn PJ=0.00041 m=1 $X=7804760 $Y=80300 $D=9
D1786 CS2 vdd! dn PJ=0.0001 m=1 $X=7805740 $Y=13228100 $D=9
D1787 CS2 vdd! dn PJ=0.0001 m=1 $X=7805740 $Y=13438100 $D=9
D1788 VDD_PAD! vdd! dn PJ=0.00041 m=1 $X=7807260 $Y=80300 $D=9
D1789 gnd! CS2 dn PJ=0.0001 m=1 $X=7808920 $Y=13332500 $D=9
D1790 gnd! CS2 dn PJ=0.0001 m=1 $X=7808920 $Y=13542500 $D=9
D1791 vdd! VDD_PAD! dn PJ=0.00041 m=1 $X=7809760 $Y=80300 $D=9
D1792 CS2 vdd! dn PJ=0.0002 m=1 $X=7811240 $Y=13228100 $D=9
D1793 CS2 vdd! dn PJ=0.0002 m=1 $X=7811240 $Y=13438100 $D=9
D1794 gnd! CS2 dn PJ=0.0002 m=1 $X=7813560 $Y=13232500 $D=9
D1795 gnd! CS2 dn PJ=0.0002 m=1 $X=7813560 $Y=13442500 $D=9
D1796 GND_PAD! VDD_PAD! dn PJ=0.00041 m=1 $X=7814760 $Y=80300 $D=9
D1797 CS2 vdd! dn PJ=0.0002 m=1 $X=7815880 $Y=13228100 $D=9
D1798 CS2 vdd! dn PJ=0.0002 m=1 $X=7815880 $Y=13438100 $D=9
D1799 VDD_PAD! vdd! dn PJ=0.00041 m=1 $X=7817260 $Y=80300 $D=9
D1800 gnd! CS2 dn PJ=0.0002 m=1 $X=7818200 $Y=13232500 $D=9
D1801 gnd! CS2 dn PJ=0.0002 m=1 $X=7818200 $Y=13442500 $D=9
D1802 vdd! VDD_PAD! dn PJ=0.00041 m=1 $X=7819760 $Y=80300 $D=9
D1803 CS2 vdd! dn PJ=0.0001 m=1 $X=7820520 $Y=13228100 $D=9
D1804 CS2 vdd! dn PJ=0.0001 m=1 $X=7820520 $Y=13438100 $D=9
D1805 gnd! CS2 dn PJ=0.0001 m=1 $X=7823700 $Y=13332500 $D=9
D1806 gnd! CS2 dn PJ=0.0001 m=1 $X=7823700 $Y=13542500 $D=9
D1807 GND_PAD! VDD_PAD! dn PJ=0.00041 m=1 $X=7824760 $Y=80300 $D=9
D1808 CS2 vdd! dn PJ=0.0002 m=1 $X=7826020 $Y=13228100 $D=9
D1809 CS2 vdd! dn PJ=0.0002 m=1 $X=7826020 $Y=13438100 $D=9
D1810 VDD_PAD! vdd! dn PJ=0.00041 m=1 $X=7827260 $Y=80300 $D=9
D1811 gnd! CS2 dn PJ=0.0002 m=1 $X=7828340 $Y=13232500 $D=9
D1812 gnd! CS2 dn PJ=0.0002 m=1 $X=7828340 $Y=13442500 $D=9
D1813 vdd! VDD_PAD! dn PJ=0.00041 m=1 $X=7829760 $Y=80300 $D=9
D1814 CS2 vdd! dn PJ=0.0002 m=1 $X=7830660 $Y=13228100 $D=9
D1815 CS2 vdd! dn PJ=0.0002 m=1 $X=7830660 $Y=13438100 $D=9
D1816 gnd! CS2 dn PJ=0.0002 m=1 $X=7832980 $Y=13232500 $D=9
D1817 gnd! CS2 dn PJ=0.0002 m=1 $X=7832980 $Y=13442500 $D=9
D1818 GND_PAD! VDD_PAD! dn PJ=0.00041 m=1 $X=7834760 $Y=80300 $D=9
D1819 CS2 vdd! dn PJ=0.0001 m=1 $X=7835300 $Y=13228100 $D=9
D1820 CS2 vdd! dn PJ=0.0001 m=1 $X=7835300 $Y=13438100 $D=9
D1821 VDD_PAD! vdd! dn PJ=0.00041 m=1 $X=7837260 $Y=80300 $D=9
D1822 gnd! CS2 dn PJ=0.0001 m=1 $X=7838480 $Y=13332500 $D=9
D1823 gnd! CS2 dn PJ=0.0001 m=1 $X=7838480 $Y=13542500 $D=9
D1824 vdd! VDD_PAD! dn PJ=0.00041 m=1 $X=7839760 $Y=80300 $D=9
D1825 CS2 vdd! dn PJ=0.0002 m=1 $X=7840800 $Y=13228100 $D=9
D1826 CS2 vdd! dn PJ=0.0002 m=1 $X=7840800 $Y=13438100 $D=9
D1827 gnd! CS2 dn PJ=0.0002 m=1 $X=7843120 $Y=13232500 $D=9
D1828 gnd! CS2 dn PJ=0.0002 m=1 $X=7843120 $Y=13442500 $D=9
D1829 GND_PAD! VDD_PAD! dn PJ=0.00041 m=1 $X=7844760 $Y=80300 $D=9
D1830 CS2 vdd! dn PJ=0.0002 m=1 $X=7845440 $Y=13228100 $D=9
D1831 CS2 vdd! dn PJ=0.0002 m=1 $X=7845440 $Y=13438100 $D=9
D1832 VDD_PAD! vdd! dn PJ=0.00041 m=1 $X=7847260 $Y=80300 $D=9
D1833 gnd! CS2 dn PJ=0.0002 m=1 $X=7847760 $Y=13232500 $D=9
D1834 gnd! CS2 dn PJ=0.0002 m=1 $X=7847760 $Y=13442500 $D=9
D1835 CS2 vdd! dn PJ=0.0001 m=1 $X=7850080 $Y=13228100 $D=9
D1836 CS2 vdd! dn PJ=0.0001 m=1 $X=7850080 $Y=13438100 $D=9
D1837 gnd! CS2 dn PJ=0.0001 m=1 $X=7853260 $Y=13332500 $D=9
D1838 gnd! CS2 dn PJ=0.0001 m=1 $X=7853260 $Y=13542500 $D=9
D1839 CS2 vdd! dn PJ=0.0002 m=1 $X=7855580 $Y=13228100 $D=9
D1840 CS2 vdd! dn PJ=0.0002 m=1 $X=7855580 $Y=13438100 $D=9
D1841 gnd! CS2 dn PJ=0.0002 m=1 $X=7857900 $Y=13232500 $D=9
D1842 gnd! CS2 dn PJ=0.0002 m=1 $X=7857900 $Y=13442500 $D=9
D1843 CS2 vdd! dn PJ=0.0002 m=1 $X=7860220 $Y=13228100 $D=9
D1844 CS2 vdd! dn PJ=0.0002 m=1 $X=7860220 $Y=13438100 $D=9
D1845 gnd! CS2 dn PJ=0.0002 m=1 $X=7862540 $Y=13232500 $D=9
D1846 gnd! CS2 dn PJ=0.0002 m=1 $X=7862540 $Y=13442500 $D=9
D1847 CS2 vdd! dn PJ=0.0001 m=1 $X=7864860 $Y=13228100 $D=9
D1848 CS2 vdd! dn PJ=0.0001 m=1 $X=7864860 $Y=13438100 $D=9
D1849 gnd! CS2 dn PJ=0.0001 m=1 $X=7868040 $Y=13332500 $D=9
D1850 gnd! CS2 dn PJ=0.0001 m=1 $X=7868040 $Y=13542500 $D=9
D1851 CS2 vdd! dn PJ=0.0002 m=1 $X=7870360 $Y=13228100 $D=9
D1852 CS2 vdd! dn PJ=0.0002 m=1 $X=7870360 $Y=13438100 $D=9
D1853 gnd! CS2 dn PJ=0.0002 m=1 $X=7872680 $Y=13232500 $D=9
D1854 gnd! CS2 dn PJ=0.0002 m=1 $X=7872680 $Y=13442500 $D=9
D1855 CS2 vdd! dn PJ=0.0002 m=1 $X=7875000 $Y=13228100 $D=9
D1856 CS2 vdd! dn PJ=0.0002 m=1 $X=7875000 $Y=13438100 $D=9
D1857 gnd! A21 dn PJ=0.0002 m=1 $X=8044000 $Y=13232500 $D=9
D1858 gnd! A21 dn PJ=0.0002 m=1 $X=8044000 $Y=13442500 $D=9
D1859 A21 vdd! dn PJ=0.0002 m=1 $X=8046320 $Y=13228100 $D=9
D1860 A21 vdd! dn PJ=0.0002 m=1 $X=8046320 $Y=13438100 $D=9
D1861 gnd! A21 dn PJ=0.0002 m=1 $X=8048640 $Y=13232500 $D=9
D1862 gnd! A21 dn PJ=0.0002 m=1 $X=8048640 $Y=13442500 $D=9
D1863 A21 vdd! dn PJ=0.0001 m=1 $X=8050960 $Y=13228100 $D=9
D1864 A21 vdd! dn PJ=0.0001 m=1 $X=8050960 $Y=13438100 $D=9
D1865 gnd! A21 dn PJ=0.0001 m=1 $X=8054140 $Y=13332500 $D=9
D1866 gnd! A21 dn PJ=0.0001 m=1 $X=8054140 $Y=13542500 $D=9
D1867 A21 vdd! dn PJ=0.0002 m=1 $X=8056460 $Y=13228100 $D=9
D1868 A21 vdd! dn PJ=0.0002 m=1 $X=8056460 $Y=13438100 $D=9
D1869 gnd! A21 dn PJ=0.0002 m=1 $X=8058780 $Y=13232500 $D=9
D1870 gnd! A21 dn PJ=0.0002 m=1 $X=8058780 $Y=13442500 $D=9
D1871 A21 vdd! dn PJ=0.0002 m=1 $X=8061100 $Y=13228100 $D=9
D1872 A21 vdd! dn PJ=0.0002 m=1 $X=8061100 $Y=13438100 $D=9
D1873 gnd! A21 dn PJ=0.0002 m=1 $X=8063420 $Y=13232500 $D=9
D1874 gnd! A21 dn PJ=0.0002 m=1 $X=8063420 $Y=13442500 $D=9
D1875 A21 vdd! dn PJ=0.0001 m=1 $X=8065740 $Y=13228100 $D=9
D1876 A21 vdd! dn PJ=0.0001 m=1 $X=8065740 $Y=13438100 $D=9
D1877 gnd! A21 dn PJ=0.0001 m=1 $X=8068920 $Y=13332500 $D=9
D1878 gnd! A21 dn PJ=0.0001 m=1 $X=8068920 $Y=13542500 $D=9
D1879 A21 vdd! dn PJ=0.0002 m=1 $X=8071240 $Y=13228100 $D=9
D1880 A21 vdd! dn PJ=0.0002 m=1 $X=8071240 $Y=13438100 $D=9
D1881 gnd! A21 dn PJ=0.0002 m=1 $X=8073560 $Y=13232500 $D=9
D1882 gnd! A21 dn PJ=0.0002 m=1 $X=8073560 $Y=13442500 $D=9
D1883 A21 vdd! dn PJ=0.0002 m=1 $X=8075880 $Y=13228100 $D=9
D1884 A21 vdd! dn PJ=0.0002 m=1 $X=8075880 $Y=13438100 $D=9
D1885 gnd! A21 dn PJ=0.0002 m=1 $X=8078200 $Y=13232500 $D=9
D1886 gnd! A21 dn PJ=0.0002 m=1 $X=8078200 $Y=13442500 $D=9
D1887 A21 vdd! dn PJ=0.0001 m=1 $X=8080520 $Y=13228100 $D=9
D1888 A21 vdd! dn PJ=0.0001 m=1 $X=8080520 $Y=13438100 $D=9
D1889 gnd! A21 dn PJ=0.0001 m=1 $X=8083700 $Y=13332500 $D=9
D1890 gnd! A21 dn PJ=0.0001 m=1 $X=8083700 $Y=13542500 $D=9
D1891 A21 vdd! dn PJ=0.0002 m=1 $X=8086020 $Y=13228100 $D=9
D1892 A21 vdd! dn PJ=0.0002 m=1 $X=8086020 $Y=13438100 $D=9
D1893 gnd! A21 dn PJ=0.0002 m=1 $X=8088340 $Y=13232500 $D=9
D1894 gnd! A21 dn PJ=0.0002 m=1 $X=8088340 $Y=13442500 $D=9
D1895 A21 vdd! dn PJ=0.0002 m=1 $X=8090660 $Y=13228100 $D=9
D1896 A21 vdd! dn PJ=0.0002 m=1 $X=8090660 $Y=13438100 $D=9
D1897 gnd! A21 dn PJ=0.0002 m=1 $X=8092980 $Y=13232500 $D=9
D1898 gnd! A21 dn PJ=0.0002 m=1 $X=8092980 $Y=13442500 $D=9
D1899 A21 vdd! dn PJ=0.0001 m=1 $X=8095300 $Y=13228100 $D=9
D1900 A21 vdd! dn PJ=0.0001 m=1 $X=8095300 $Y=13438100 $D=9
D1901 gnd! A21 dn PJ=0.0001 m=1 $X=8098480 $Y=13332500 $D=9
D1902 gnd! A21 dn PJ=0.0001 m=1 $X=8098480 $Y=13542500 $D=9
D1903 A21 vdd! dn PJ=0.0002 m=1 $X=8100800 $Y=13228100 $D=9
D1904 A21 vdd! dn PJ=0.0002 m=1 $X=8100800 $Y=13438100 $D=9
D1905 gnd! A21 dn PJ=0.0002 m=1 $X=8103120 $Y=13232500 $D=9
D1906 gnd! A21 dn PJ=0.0002 m=1 $X=8103120 $Y=13442500 $D=9
D1907 A21 vdd! dn PJ=0.0002 m=1 $X=8105440 $Y=13228100 $D=9
D1908 A21 vdd! dn PJ=0.0002 m=1 $X=8105440 $Y=13438100 $D=9
D1909 gnd! A21 dn PJ=0.0002 m=1 $X=8107760 $Y=13232500 $D=9
D1910 gnd! A21 dn PJ=0.0002 m=1 $X=8107760 $Y=13442500 $D=9
D1911 A21 vdd! dn PJ=0.0001 m=1 $X=8110080 $Y=13228100 $D=9
D1912 A21 vdd! dn PJ=0.0001 m=1 $X=8110080 $Y=13438100 $D=9
D1913 gnd! A21 dn PJ=0.0001 m=1 $X=8113260 $Y=13332500 $D=9
D1914 gnd! A21 dn PJ=0.0001 m=1 $X=8113260 $Y=13542500 $D=9
D1915 A21 vdd! dn PJ=0.0002 m=1 $X=8115580 $Y=13228100 $D=9
D1916 A21 vdd! dn PJ=0.0002 m=1 $X=8115580 $Y=13438100 $D=9
D1917 gnd! A21 dn PJ=0.0002 m=1 $X=8117900 $Y=13232500 $D=9
D1918 gnd! A21 dn PJ=0.0002 m=1 $X=8117900 $Y=13442500 $D=9
D1919 A21 vdd! dn PJ=0.0002 m=1 $X=8120220 $Y=13228100 $D=9
D1920 A21 vdd! dn PJ=0.0002 m=1 $X=8120220 $Y=13438100 $D=9
D1921 gnd! A21 dn PJ=0.0002 m=1 $X=8122540 $Y=13232500 $D=9
D1922 gnd! A21 dn PJ=0.0002 m=1 $X=8122540 $Y=13442500 $D=9
D1923 A21 vdd! dn PJ=0.0001 m=1 $X=8124860 $Y=13228100 $D=9
D1924 A21 vdd! dn PJ=0.0001 m=1 $X=8124860 $Y=13438100 $D=9
D1925 gnd! A21 dn PJ=0.0001 m=1 $X=8128040 $Y=13332500 $D=9
D1926 gnd! A21 dn PJ=0.0001 m=1 $X=8128040 $Y=13542500 $D=9
D1927 A21 vdd! dn PJ=0.0002 m=1 $X=8130360 $Y=13228100 $D=9
D1928 A21 vdd! dn PJ=0.0002 m=1 $X=8130360 $Y=13438100 $D=9
D1929 gnd! A21 dn PJ=0.0002 m=1 $X=8132680 $Y=13232500 $D=9
D1930 gnd! A21 dn PJ=0.0002 m=1 $X=8132680 $Y=13442500 $D=9
D1931 A21 vdd! dn PJ=0.0002 m=1 $X=8135000 $Y=13228100 $D=9
D1932 A21 vdd! dn PJ=0.0002 m=1 $X=8135000 $Y=13438100 $D=9
D1933 gnd! A12 dn PJ=0.0002 m=1 $X=10124000 $Y=13232500 $D=9
D1934 gnd! A12 dn PJ=0.0002 m=1 $X=10124000 $Y=13442500 $D=9
D1935 A12 vdd! dn PJ=0.0002 m=1 $X=10126320 $Y=13228100 $D=9
D1936 A12 vdd! dn PJ=0.0002 m=1 $X=10126320 $Y=13438100 $D=9
D1937 gnd! A12 dn PJ=0.0002 m=1 $X=10128640 $Y=13232500 $D=9
D1938 gnd! A12 dn PJ=0.0002 m=1 $X=10128640 $Y=13442500 $D=9
D1939 A12 vdd! dn PJ=0.0001 m=1 $X=10130960 $Y=13228100 $D=9
D1940 A12 vdd! dn PJ=0.0001 m=1 $X=10130960 $Y=13438100 $D=9
D1941 gnd! A12 dn PJ=0.0001 m=1 $X=10134140 $Y=13332500 $D=9
D1942 gnd! A12 dn PJ=0.0001 m=1 $X=10134140 $Y=13542500 $D=9
D1943 A12 vdd! dn PJ=0.0002 m=1 $X=10136460 $Y=13228100 $D=9
D1944 A12 vdd! dn PJ=0.0002 m=1 $X=10136460 $Y=13438100 $D=9
D1945 gnd! A12 dn PJ=0.0002 m=1 $X=10138780 $Y=13232500 $D=9
D1946 gnd! A12 dn PJ=0.0002 m=1 $X=10138780 $Y=13442500 $D=9
D1947 A12 vdd! dn PJ=0.0002 m=1 $X=10141100 $Y=13228100 $D=9
D1948 A12 vdd! dn PJ=0.0002 m=1 $X=10141100 $Y=13438100 $D=9
D1949 gnd! A12 dn PJ=0.0002 m=1 $X=10143420 $Y=13232500 $D=9
D1950 gnd! A12 dn PJ=0.0002 m=1 $X=10143420 $Y=13442500 $D=9
D1951 A12 vdd! dn PJ=0.0001 m=1 $X=10145740 $Y=13228100 $D=9
D1952 A12 vdd! dn PJ=0.0001 m=1 $X=10145740 $Y=13438100 $D=9
D1953 gnd! A12 dn PJ=0.0001 m=1 $X=10148920 $Y=13332500 $D=9
D1954 gnd! A12 dn PJ=0.0001 m=1 $X=10148920 $Y=13542500 $D=9
D1955 A12 vdd! dn PJ=0.0002 m=1 $X=10151240 $Y=13228100 $D=9
D1956 A12 vdd! dn PJ=0.0002 m=1 $X=10151240 $Y=13438100 $D=9
D1957 gnd! A12 dn PJ=0.0002 m=1 $X=10153560 $Y=13232500 $D=9
D1958 gnd! A12 dn PJ=0.0002 m=1 $X=10153560 $Y=13442500 $D=9
D1959 A12 vdd! dn PJ=0.0002 m=1 $X=10155880 $Y=13228100 $D=9
D1960 A12 vdd! dn PJ=0.0002 m=1 $X=10155880 $Y=13438100 $D=9
D1961 gnd! A12 dn PJ=0.0002 m=1 $X=10158200 $Y=13232500 $D=9
D1962 gnd! A12 dn PJ=0.0002 m=1 $X=10158200 $Y=13442500 $D=9
D1963 A12 vdd! dn PJ=0.0001 m=1 $X=10160520 $Y=13228100 $D=9
D1964 A12 vdd! dn PJ=0.0001 m=1 $X=10160520 $Y=13438100 $D=9
D1965 gnd! A12 dn PJ=0.0001 m=1 $X=10163700 $Y=13332500 $D=9
D1966 gnd! A12 dn PJ=0.0001 m=1 $X=10163700 $Y=13542500 $D=9
D1967 A12 vdd! dn PJ=0.0002 m=1 $X=10166020 $Y=13228100 $D=9
D1968 A12 vdd! dn PJ=0.0002 m=1 $X=10166020 $Y=13438100 $D=9
D1969 gnd! A12 dn PJ=0.0002 m=1 $X=10168340 $Y=13232500 $D=9
D1970 gnd! A12 dn PJ=0.0002 m=1 $X=10168340 $Y=13442500 $D=9
D1971 A12 vdd! dn PJ=0.0002 m=1 $X=10170660 $Y=13228100 $D=9
D1972 A12 vdd! dn PJ=0.0002 m=1 $X=10170660 $Y=13438100 $D=9
D1973 gnd! A12 dn PJ=0.0002 m=1 $X=10172980 $Y=13232500 $D=9
D1974 gnd! A12 dn PJ=0.0002 m=1 $X=10172980 $Y=13442500 $D=9
D1975 A12 vdd! dn PJ=0.0001 m=1 $X=10175300 $Y=13228100 $D=9
D1976 A12 vdd! dn PJ=0.0001 m=1 $X=10175300 $Y=13438100 $D=9
D1977 gnd! A12 dn PJ=0.0001 m=1 $X=10178480 $Y=13332500 $D=9
D1978 gnd! A12 dn PJ=0.0001 m=1 $X=10178480 $Y=13542500 $D=9
D1979 A12 vdd! dn PJ=0.0002 m=1 $X=10180800 $Y=13228100 $D=9
D1980 A12 vdd! dn PJ=0.0002 m=1 $X=10180800 $Y=13438100 $D=9
D1981 gnd! A12 dn PJ=0.0002 m=1 $X=10183120 $Y=13232500 $D=9
D1982 gnd! A12 dn PJ=0.0002 m=1 $X=10183120 $Y=13442500 $D=9
D1983 A12 vdd! dn PJ=0.0002 m=1 $X=10185440 $Y=13228100 $D=9
D1984 A12 vdd! dn PJ=0.0002 m=1 $X=10185440 $Y=13438100 $D=9
D1985 gnd! A12 dn PJ=0.0002 m=1 $X=10187760 $Y=13232500 $D=9
D1986 gnd! A12 dn PJ=0.0002 m=1 $X=10187760 $Y=13442500 $D=9
D1987 A12 vdd! dn PJ=0.0001 m=1 $X=10190080 $Y=13228100 $D=9
D1988 A12 vdd! dn PJ=0.0001 m=1 $X=10190080 $Y=13438100 $D=9
D1989 gnd! A12 dn PJ=0.0001 m=1 $X=10193260 $Y=13332500 $D=9
D1990 gnd! A12 dn PJ=0.0001 m=1 $X=10193260 $Y=13542500 $D=9
D1991 A12 vdd! dn PJ=0.0002 m=1 $X=10195580 $Y=13228100 $D=9
D1992 A12 vdd! dn PJ=0.0002 m=1 $X=10195580 $Y=13438100 $D=9
D1993 gnd! A12 dn PJ=0.0002 m=1 $X=10197900 $Y=13232500 $D=9
D1994 gnd! A12 dn PJ=0.0002 m=1 $X=10197900 $Y=13442500 $D=9
D1995 A12 vdd! dn PJ=0.0002 m=1 $X=10200220 $Y=13228100 $D=9
D1996 A12 vdd! dn PJ=0.0002 m=1 $X=10200220 $Y=13438100 $D=9
D1997 gnd! A12 dn PJ=0.0002 m=1 $X=10202540 $Y=13232500 $D=9
D1998 gnd! A12 dn PJ=0.0002 m=1 $X=10202540 $Y=13442500 $D=9
D1999 A12 vdd! dn PJ=0.0001 m=1 $X=10204860 $Y=13228100 $D=9
D2000 A12 vdd! dn PJ=0.0001 m=1 $X=10204860 $Y=13438100 $D=9
D2001 gnd! A12 dn PJ=0.0001 m=1 $X=10208040 $Y=13332500 $D=9
D2002 gnd! A12 dn PJ=0.0001 m=1 $X=10208040 $Y=13542500 $D=9
D2003 A12 vdd! dn PJ=0.0002 m=1 $X=10210360 $Y=13228100 $D=9
D2004 A12 vdd! dn PJ=0.0002 m=1 $X=10210360 $Y=13438100 $D=9
D2005 gnd! A12 dn PJ=0.0002 m=1 $X=10212680 $Y=13232500 $D=9
D2006 gnd! A12 dn PJ=0.0002 m=1 $X=10212680 $Y=13442500 $D=9
D2007 A12 vdd! dn PJ=0.0002 m=1 $X=10215000 $Y=13228100 $D=9
D2008 A12 vdd! dn PJ=0.0002 m=1 $X=10215000 $Y=13438100 $D=9
D2009 GND_PAD! VDD_PAD! dn PJ=0.00041 m=1 $X=10454760 $Y=80300 $D=9
D2010 VDD_PAD! vdd! dn PJ=0.00041 m=1 $X=10457260 $Y=80300 $D=9
D2011 vdd! VDD_PAD! dn PJ=0.00041 m=1 $X=10459760 $Y=80300 $D=9
D2012 GND_PAD! VDD_PAD! dn PJ=0.00041 m=1 $X=10464760 $Y=80300 $D=9
D2013 VDD_PAD! vdd! dn PJ=0.00041 m=1 $X=10467260 $Y=80300 $D=9
D2014 vdd! VDD_PAD! dn PJ=0.00041 m=1 $X=10469760 $Y=80300 $D=9
D2015 GND_PAD! VDD_PAD! dn PJ=0.00041 m=1 $X=10474760 $Y=80300 $D=9
D2016 VDD_PAD! vdd! dn PJ=0.00041 m=1 $X=10477260 $Y=80300 $D=9
D2017 vdd! VDD_PAD! dn PJ=0.00041 m=1 $X=10479760 $Y=80300 $D=9
D2018 GND_PAD! VDD_PAD! dn PJ=0.00041 m=1 $X=10484760 $Y=80300 $D=9
D2019 VDD_PAD! vdd! dn PJ=0.00041 m=1 $X=10487260 $Y=80300 $D=9
D2020 vdd! VDD_PAD! dn PJ=0.00041 m=1 $X=10489760 $Y=80300 $D=9
D2021 GND_PAD! VDD_PAD! dn PJ=0.00041 m=1 $X=10494760 $Y=80300 $D=9
D2022 VDD_PAD! vdd! dn PJ=0.00041 m=1 $X=10497260 $Y=80300 $D=9
D2023 vdd! VDD_PAD! dn PJ=0.00041 m=1 $X=10499760 $Y=80300 $D=9
D2024 GND_PAD! VDD_PAD! dn PJ=0.00041 m=1 $X=10504760 $Y=80300 $D=9
D2025 VDD_PAD! vdd! dn PJ=0.00041 m=1 $X=10507260 $Y=80300 $D=9
D2026 vdd! VDD_PAD! dn PJ=0.00041 m=1 $X=10509760 $Y=80300 $D=9
D2027 GND_PAD! VDD_PAD! dn PJ=0.00041 m=1 $X=10514760 $Y=80300 $D=9
D2028 VDD_PAD! vdd! dn PJ=0.00041 m=1 $X=10517260 $Y=80300 $D=9
D2029 vdd! VDD_PAD! dn PJ=0.00041 m=1 $X=10519760 $Y=80300 $D=9
D2030 GND_PAD! VDD_PAD! dn PJ=0.00041 m=1 $X=10524760 $Y=80300 $D=9
D2031 VDD_PAD! vdd! dn PJ=0.00041 m=1 $X=10527260 $Y=80300 $D=9
D2032 vdd! VDD_PAD! dn PJ=0.00041 m=1 $X=10529760 $Y=80300 $D=9
D2033 GND_PAD! VDD_PAD! dn PJ=0.00041 m=1 $X=10534760 $Y=80300 $D=9
D2034 VDD_PAD! vdd! dn PJ=0.00041 m=1 $X=10537260 $Y=80300 $D=9
D2035 vdd! VDD_PAD! dn PJ=0.00041 m=1 $X=10539760 $Y=80300 $D=9
D2036 GND_PAD! VDD_PAD! dn PJ=0.00041 m=1 $X=10544760 $Y=80300 $D=9
D2037 VDD_PAD! vdd! dn PJ=0.00041 m=1 $X=10547260 $Y=80300 $D=9
D2038 gnd! A14 dn PJ=0.0002 m=1 $X=10644000 $Y=13232500 $D=9
D2039 gnd! A14 dn PJ=0.0002 m=1 $X=10644000 $Y=13442500 $D=9
D2040 A14 vdd! dn PJ=0.0002 m=1 $X=10646320 $Y=13228100 $D=9
D2041 A14 vdd! dn PJ=0.0002 m=1 $X=10646320 $Y=13438100 $D=9
D2042 gnd! A14 dn PJ=0.0002 m=1 $X=10648640 $Y=13232500 $D=9
D2043 gnd! A14 dn PJ=0.0002 m=1 $X=10648640 $Y=13442500 $D=9
D2044 A14 vdd! dn PJ=0.0001 m=1 $X=10650960 $Y=13228100 $D=9
D2045 A14 vdd! dn PJ=0.0001 m=1 $X=10650960 $Y=13438100 $D=9
D2046 gnd! A14 dn PJ=0.0001 m=1 $X=10654140 $Y=13332500 $D=9
D2047 gnd! A14 dn PJ=0.0001 m=1 $X=10654140 $Y=13542500 $D=9
D2048 A14 vdd! dn PJ=0.0002 m=1 $X=10656460 $Y=13228100 $D=9
D2049 A14 vdd! dn PJ=0.0002 m=1 $X=10656460 $Y=13438100 $D=9
D2050 gnd! A14 dn PJ=0.0002 m=1 $X=10658780 $Y=13232500 $D=9
D2051 gnd! A14 dn PJ=0.0002 m=1 $X=10658780 $Y=13442500 $D=9
D2052 A14 vdd! dn PJ=0.0002 m=1 $X=10661100 $Y=13228100 $D=9
D2053 A14 vdd! dn PJ=0.0002 m=1 $X=10661100 $Y=13438100 $D=9
D2054 gnd! A14 dn PJ=0.0002 m=1 $X=10663420 $Y=13232500 $D=9
D2055 gnd! A14 dn PJ=0.0002 m=1 $X=10663420 $Y=13442500 $D=9
D2056 A14 vdd! dn PJ=0.0001 m=1 $X=10665740 $Y=13228100 $D=9
D2057 A14 vdd! dn PJ=0.0001 m=1 $X=10665740 $Y=13438100 $D=9
D2058 gnd! A14 dn PJ=0.0001 m=1 $X=10668920 $Y=13332500 $D=9
D2059 gnd! A14 dn PJ=0.0001 m=1 $X=10668920 $Y=13542500 $D=9
D2060 A14 vdd! dn PJ=0.0002 m=1 $X=10671240 $Y=13228100 $D=9
D2061 A14 vdd! dn PJ=0.0002 m=1 $X=10671240 $Y=13438100 $D=9
D2062 gnd! A14 dn PJ=0.0002 m=1 $X=10673560 $Y=13232500 $D=9
D2063 gnd! A14 dn PJ=0.0002 m=1 $X=10673560 $Y=13442500 $D=9
D2064 A14 vdd! dn PJ=0.0002 m=1 $X=10675880 $Y=13228100 $D=9
D2065 A14 vdd! dn PJ=0.0002 m=1 $X=10675880 $Y=13438100 $D=9
D2066 gnd! A14 dn PJ=0.0002 m=1 $X=10678200 $Y=13232500 $D=9
D2067 gnd! A14 dn PJ=0.0002 m=1 $X=10678200 $Y=13442500 $D=9
D2068 A14 vdd! dn PJ=0.0001 m=1 $X=10680520 $Y=13228100 $D=9
D2069 A14 vdd! dn PJ=0.0001 m=1 $X=10680520 $Y=13438100 $D=9
D2070 gnd! A14 dn PJ=0.0001 m=1 $X=10683700 $Y=13332500 $D=9
D2071 gnd! A14 dn PJ=0.0001 m=1 $X=10683700 $Y=13542500 $D=9
D2072 A14 vdd! dn PJ=0.0002 m=1 $X=10686020 $Y=13228100 $D=9
D2073 A14 vdd! dn PJ=0.0002 m=1 $X=10686020 $Y=13438100 $D=9
D2074 gnd! A14 dn PJ=0.0002 m=1 $X=10688340 $Y=13232500 $D=9
D2075 gnd! A14 dn PJ=0.0002 m=1 $X=10688340 $Y=13442500 $D=9
D2076 A14 vdd! dn PJ=0.0002 m=1 $X=10690660 $Y=13228100 $D=9
D2077 A14 vdd! dn PJ=0.0002 m=1 $X=10690660 $Y=13438100 $D=9
D2078 gnd! A14 dn PJ=0.0002 m=1 $X=10692980 $Y=13232500 $D=9
D2079 gnd! A14 dn PJ=0.0002 m=1 $X=10692980 $Y=13442500 $D=9
D2080 A14 vdd! dn PJ=0.0001 m=1 $X=10695300 $Y=13228100 $D=9
D2081 A14 vdd! dn PJ=0.0001 m=1 $X=10695300 $Y=13438100 $D=9
D2082 gnd! A14 dn PJ=0.0001 m=1 $X=10698480 $Y=13332500 $D=9
D2083 gnd! A14 dn PJ=0.0001 m=1 $X=10698480 $Y=13542500 $D=9
D2084 A14 vdd! dn PJ=0.0002 m=1 $X=10700800 $Y=13228100 $D=9
D2085 A14 vdd! dn PJ=0.0002 m=1 $X=10700800 $Y=13438100 $D=9
D2086 gnd! A14 dn PJ=0.0002 m=1 $X=10703120 $Y=13232500 $D=9
D2087 gnd! A14 dn PJ=0.0002 m=1 $X=10703120 $Y=13442500 $D=9
D2088 A14 vdd! dn PJ=0.0002 m=1 $X=10705440 $Y=13228100 $D=9
D2089 A14 vdd! dn PJ=0.0002 m=1 $X=10705440 $Y=13438100 $D=9
D2090 gnd! A14 dn PJ=0.0002 m=1 $X=10707760 $Y=13232500 $D=9
D2091 gnd! A14 dn PJ=0.0002 m=1 $X=10707760 $Y=13442500 $D=9
D2092 A14 vdd! dn PJ=0.0001 m=1 $X=10710080 $Y=13228100 $D=9
D2093 A14 vdd! dn PJ=0.0001 m=1 $X=10710080 $Y=13438100 $D=9
D2094 gnd! A14 dn PJ=0.0001 m=1 $X=10713260 $Y=13332500 $D=9
D2095 gnd! A14 dn PJ=0.0001 m=1 $X=10713260 $Y=13542500 $D=9
D2096 A14 vdd! dn PJ=0.0002 m=1 $X=10715580 $Y=13228100 $D=9
D2097 A14 vdd! dn PJ=0.0002 m=1 $X=10715580 $Y=13438100 $D=9
D2098 gnd! A14 dn PJ=0.0002 m=1 $X=10717900 $Y=13232500 $D=9
D2099 gnd! A14 dn PJ=0.0002 m=1 $X=10717900 $Y=13442500 $D=9
D2100 A14 vdd! dn PJ=0.0002 m=1 $X=10720220 $Y=13228100 $D=9
D2101 A14 vdd! dn PJ=0.0002 m=1 $X=10720220 $Y=13438100 $D=9
D2102 gnd! A14 dn PJ=0.0002 m=1 $X=10722540 $Y=13232500 $D=9
D2103 gnd! A14 dn PJ=0.0002 m=1 $X=10722540 $Y=13442500 $D=9
D2104 A14 vdd! dn PJ=0.0001 m=1 $X=10724860 $Y=13228100 $D=9
D2105 A14 vdd! dn PJ=0.0001 m=1 $X=10724860 $Y=13438100 $D=9
D2106 gnd! A14 dn PJ=0.0001 m=1 $X=10728040 $Y=13332500 $D=9
D2107 gnd! A14 dn PJ=0.0001 m=1 $X=10728040 $Y=13542500 $D=9
D2108 A14 vdd! dn PJ=0.0002 m=1 $X=10730360 $Y=13228100 $D=9
D2109 A14 vdd! dn PJ=0.0002 m=1 $X=10730360 $Y=13438100 $D=9
D2110 gnd! A14 dn PJ=0.0002 m=1 $X=10732680 $Y=13232500 $D=9
D2111 gnd! A14 dn PJ=0.0002 m=1 $X=10732680 $Y=13442500 $D=9
D2112 A14 vdd! dn PJ=0.0002 m=1 $X=10735000 $Y=13228100 $D=9
D2113 A14 vdd! dn PJ=0.0002 m=1 $X=10735000 $Y=13438100 $D=9
D2114 GND_PAD! VDD_PAD! dn PJ=0.00041 m=1 $X=10754760 $Y=80300 $D=9
D2115 VDD_PAD! vdd! dn PJ=0.00041 m=1 $X=10757260 $Y=80300 $D=9
D2116 vdd! VDD_PAD! dn PJ=0.00041 m=1 $X=10759760 $Y=80300 $D=9
D2117 GND_PAD! VDD_PAD! dn PJ=0.00041 m=1 $X=10764760 $Y=80300 $D=9
D2118 VDD_PAD! vdd! dn PJ=0.00041 m=1 $X=10767260 $Y=80300 $D=9
D2119 vdd! VDD_PAD! dn PJ=0.00041 m=1 $X=10769760 $Y=80300 $D=9
D2120 GND_PAD! VDD_PAD! dn PJ=0.00041 m=1 $X=10774760 $Y=80300 $D=9
D2121 VDD_PAD! vdd! dn PJ=0.00041 m=1 $X=10777260 $Y=80300 $D=9
D2122 vdd! VDD_PAD! dn PJ=0.00041 m=1 $X=10779760 $Y=80300 $D=9
D2123 GND_PAD! VDD_PAD! dn PJ=0.00041 m=1 $X=10784760 $Y=80300 $D=9
D2124 VDD_PAD! vdd! dn PJ=0.00041 m=1 $X=10787260 $Y=80300 $D=9
D2125 vdd! VDD_PAD! dn PJ=0.00041 m=1 $X=10789760 $Y=80300 $D=9
D2126 GND_PAD! VDD_PAD! dn PJ=0.00041 m=1 $X=10794760 $Y=80300 $D=9
D2127 VDD_PAD! vdd! dn PJ=0.00041 m=1 $X=10797260 $Y=80300 $D=9
D2128 vdd! VDD_PAD! dn PJ=0.00041 m=1 $X=10799760 $Y=80300 $D=9
D2129 GND_PAD! VDD_PAD! dn PJ=0.00041 m=1 $X=10804760 $Y=80300 $D=9
D2130 VDD_PAD! vdd! dn PJ=0.00041 m=1 $X=10807260 $Y=80300 $D=9
D2131 vdd! VDD_PAD! dn PJ=0.00041 m=1 $X=10809760 $Y=80300 $D=9
D2132 GND_PAD! VDD_PAD! dn PJ=0.00041 m=1 $X=10814760 $Y=80300 $D=9
D2133 VDD_PAD! vdd! dn PJ=0.00041 m=1 $X=10817260 $Y=80300 $D=9
D2134 vdd! VDD_PAD! dn PJ=0.00041 m=1 $X=10819760 $Y=80300 $D=9
D2135 GND_PAD! VDD_PAD! dn PJ=0.00041 m=1 $X=10824760 $Y=80300 $D=9
D2136 VDD_PAD! vdd! dn PJ=0.00041 m=1 $X=10827260 $Y=80300 $D=9
D2137 vdd! VDD_PAD! dn PJ=0.00041 m=1 $X=10829760 $Y=80300 $D=9
D2138 GND_PAD! VDD_PAD! dn PJ=0.00041 m=1 $X=10834760 $Y=80300 $D=9
D2139 VDD_PAD! vdd! dn PJ=0.00041 m=1 $X=10837260 $Y=80300 $D=9
D2140 vdd! VDD_PAD! dn PJ=0.00041 m=1 $X=10839760 $Y=80300 $D=9
D2141 GND_PAD! VDD_PAD! dn PJ=0.00041 m=1 $X=10844760 $Y=80300 $D=9
D2142 VDD_PAD! vdd! dn PJ=0.00041 m=1 $X=10847260 $Y=80300 $D=9
D2143 gnd! A17 dn PJ=0.0002 m=1 $X=11944000 $Y=13232500 $D=9
D2144 gnd! A17 dn PJ=0.0002 m=1 $X=11944000 $Y=13442500 $D=9
D2145 A17 vdd! dn PJ=0.0002 m=1 $X=11946320 $Y=13228100 $D=9
D2146 A17 vdd! dn PJ=0.0002 m=1 $X=11946320 $Y=13438100 $D=9
D2147 gnd! A17 dn PJ=0.0002 m=1 $X=11948640 $Y=13232500 $D=9
D2148 gnd! A17 dn PJ=0.0002 m=1 $X=11948640 $Y=13442500 $D=9
D2149 A17 vdd! dn PJ=0.0001 m=1 $X=11950960 $Y=13228100 $D=9
D2150 A17 vdd! dn PJ=0.0001 m=1 $X=11950960 $Y=13438100 $D=9
D2151 gnd! A17 dn PJ=0.0001 m=1 $X=11954140 $Y=13332500 $D=9
D2152 gnd! A17 dn PJ=0.0001 m=1 $X=11954140 $Y=13542500 $D=9
D2153 A17 vdd! dn PJ=0.0002 m=1 $X=11956460 $Y=13228100 $D=9
D2154 A17 vdd! dn PJ=0.0002 m=1 $X=11956460 $Y=13438100 $D=9
D2155 gnd! A17 dn PJ=0.0002 m=1 $X=11958780 $Y=13232500 $D=9
D2156 gnd! A17 dn PJ=0.0002 m=1 $X=11958780 $Y=13442500 $D=9
D2157 A17 vdd! dn PJ=0.0002 m=1 $X=11961100 $Y=13228100 $D=9
D2158 A17 vdd! dn PJ=0.0002 m=1 $X=11961100 $Y=13438100 $D=9
D2159 gnd! A17 dn PJ=0.0002 m=1 $X=11963420 $Y=13232500 $D=9
D2160 gnd! A17 dn PJ=0.0002 m=1 $X=11963420 $Y=13442500 $D=9
D2161 A17 vdd! dn PJ=0.0001 m=1 $X=11965740 $Y=13228100 $D=9
D2162 A17 vdd! dn PJ=0.0001 m=1 $X=11965740 $Y=13438100 $D=9
D2163 gnd! A17 dn PJ=0.0001 m=1 $X=11968920 $Y=13332500 $D=9
D2164 gnd! A17 dn PJ=0.0001 m=1 $X=11968920 $Y=13542500 $D=9
D2165 A17 vdd! dn PJ=0.0002 m=1 $X=11971240 $Y=13228100 $D=9
D2166 A17 vdd! dn PJ=0.0002 m=1 $X=11971240 $Y=13438100 $D=9
D2167 gnd! A17 dn PJ=0.0002 m=1 $X=11973560 $Y=13232500 $D=9
D2168 gnd! A17 dn PJ=0.0002 m=1 $X=11973560 $Y=13442500 $D=9
D2169 A17 vdd! dn PJ=0.0002 m=1 $X=11975880 $Y=13228100 $D=9
D2170 A17 vdd! dn PJ=0.0002 m=1 $X=11975880 $Y=13438100 $D=9
D2171 gnd! A17 dn PJ=0.0002 m=1 $X=11978200 $Y=13232500 $D=9
D2172 gnd! A17 dn PJ=0.0002 m=1 $X=11978200 $Y=13442500 $D=9
D2173 A17 vdd! dn PJ=0.0001 m=1 $X=11980520 $Y=13228100 $D=9
D2174 A17 vdd! dn PJ=0.0001 m=1 $X=11980520 $Y=13438100 $D=9
D2175 gnd! A17 dn PJ=0.0001 m=1 $X=11983700 $Y=13332500 $D=9
D2176 gnd! A17 dn PJ=0.0001 m=1 $X=11983700 $Y=13542500 $D=9
D2177 A17 vdd! dn PJ=0.0002 m=1 $X=11986020 $Y=13228100 $D=9
D2178 A17 vdd! dn PJ=0.0002 m=1 $X=11986020 $Y=13438100 $D=9
D2179 gnd! A17 dn PJ=0.0002 m=1 $X=11988340 $Y=13232500 $D=9
D2180 gnd! A17 dn PJ=0.0002 m=1 $X=11988340 $Y=13442500 $D=9
D2181 A17 vdd! dn PJ=0.0002 m=1 $X=11990660 $Y=13228100 $D=9
D2182 A17 vdd! dn PJ=0.0002 m=1 $X=11990660 $Y=13438100 $D=9
D2183 gnd! A17 dn PJ=0.0002 m=1 $X=11992980 $Y=13232500 $D=9
D2184 gnd! A17 dn PJ=0.0002 m=1 $X=11992980 $Y=13442500 $D=9
D2185 A17 vdd! dn PJ=0.0001 m=1 $X=11995300 $Y=13228100 $D=9
D2186 A17 vdd! dn PJ=0.0001 m=1 $X=11995300 $Y=13438100 $D=9
D2187 gnd! A17 dn PJ=0.0001 m=1 $X=11998480 $Y=13332500 $D=9
D2188 gnd! A17 dn PJ=0.0001 m=1 $X=11998480 $Y=13542500 $D=9
D2189 A17 vdd! dn PJ=0.0002 m=1 $X=12000800 $Y=13228100 $D=9
D2190 A17 vdd! dn PJ=0.0002 m=1 $X=12000800 $Y=13438100 $D=9
D2191 gnd! A17 dn PJ=0.0002 m=1 $X=12003120 $Y=13232500 $D=9
D2192 gnd! A17 dn PJ=0.0002 m=1 $X=12003120 $Y=13442500 $D=9
D2193 A17 vdd! dn PJ=0.0002 m=1 $X=12005440 $Y=13228100 $D=9
D2194 A17 vdd! dn PJ=0.0002 m=1 $X=12005440 $Y=13438100 $D=9
D2195 gnd! A17 dn PJ=0.0002 m=1 $X=12007760 $Y=13232500 $D=9
D2196 gnd! A17 dn PJ=0.0002 m=1 $X=12007760 $Y=13442500 $D=9
D2197 A17 vdd! dn PJ=0.0001 m=1 $X=12010080 $Y=13228100 $D=9
D2198 A17 vdd! dn PJ=0.0001 m=1 $X=12010080 $Y=13438100 $D=9
D2199 gnd! A17 dn PJ=0.0001 m=1 $X=12013260 $Y=13332500 $D=9
D2200 gnd! A17 dn PJ=0.0001 m=1 $X=12013260 $Y=13542500 $D=9
D2201 A17 vdd! dn PJ=0.0002 m=1 $X=12015580 $Y=13228100 $D=9
D2202 A17 vdd! dn PJ=0.0002 m=1 $X=12015580 $Y=13438100 $D=9
D2203 gnd! A17 dn PJ=0.0002 m=1 $X=12017900 $Y=13232500 $D=9
D2204 gnd! A17 dn PJ=0.0002 m=1 $X=12017900 $Y=13442500 $D=9
D2205 A17 vdd! dn PJ=0.0002 m=1 $X=12020220 $Y=13228100 $D=9
D2206 A17 vdd! dn PJ=0.0002 m=1 $X=12020220 $Y=13438100 $D=9
D2207 gnd! A17 dn PJ=0.0002 m=1 $X=12022540 $Y=13232500 $D=9
D2208 gnd! A17 dn PJ=0.0002 m=1 $X=12022540 $Y=13442500 $D=9
D2209 A17 vdd! dn PJ=0.0001 m=1 $X=12024860 $Y=13228100 $D=9
D2210 A17 vdd! dn PJ=0.0001 m=1 $X=12024860 $Y=13438100 $D=9
D2211 gnd! A17 dn PJ=0.0001 m=1 $X=12028040 $Y=13332500 $D=9
D2212 gnd! A17 dn PJ=0.0001 m=1 $X=12028040 $Y=13542500 $D=9
D2213 A17 vdd! dn PJ=0.0002 m=1 $X=12030360 $Y=13228100 $D=9
D2214 A17 vdd! dn PJ=0.0002 m=1 $X=12030360 $Y=13438100 $D=9
D2215 gnd! A17 dn PJ=0.0002 m=1 $X=12032680 $Y=13232500 $D=9
D2216 gnd! A17 dn PJ=0.0002 m=1 $X=12032680 $Y=13442500 $D=9
D2217 A17 vdd! dn PJ=0.0002 m=1 $X=12035000 $Y=13228100 $D=9
D2218 A17 vdd! dn PJ=0.0002 m=1 $X=12035000 $Y=13438100 $D=9
D2219 GND_PAD! VDD_PAD! dn PJ=0.00041 m=1 $X=14054760 $Y=80300 $D=9
D2220 VDD_PAD! vdd! dn PJ=0.00041 m=1 $X=14057260 $Y=80300 $D=9
D2221 vdd! VDD_PAD! dn PJ=0.00041 m=1 $X=14059760 $Y=80300 $D=9
D2222 GND_PAD! VDD_PAD! dn PJ=0.00041 m=1 $X=14064760 $Y=80300 $D=9
D2223 VDD_PAD! vdd! dn PJ=0.00041 m=1 $X=14067260 $Y=80300 $D=9
D2224 vdd! VDD_PAD! dn PJ=0.00041 m=1 $X=14069760 $Y=80300 $D=9
D2225 GND_PAD! VDD_PAD! dn PJ=0.00041 m=1 $X=14074760 $Y=80300 $D=9
D2226 VDD_PAD! vdd! dn PJ=0.00041 m=1 $X=14077260 $Y=80300 $D=9
D2227 vdd! VDD_PAD! dn PJ=0.00041 m=1 $X=14079760 $Y=80300 $D=9
D2228 GND_PAD! VDD_PAD! dn PJ=0.00041 m=1 $X=14084760 $Y=80300 $D=9
D2229 VDD_PAD! vdd! dn PJ=0.00041 m=1 $X=14087260 $Y=80300 $D=9
D2230 vdd! VDD_PAD! dn PJ=0.00041 m=1 $X=14089760 $Y=80300 $D=9
D2231 GND_PAD! VDD_PAD! dn PJ=0.00041 m=1 $X=14094760 $Y=80300 $D=9
D2232 VDD_PAD! vdd! dn PJ=0.00041 m=1 $X=14097260 $Y=80300 $D=9
D2233 vdd! VDD_PAD! dn PJ=0.00041 m=1 $X=14099760 $Y=80300 $D=9
D2234 GND_PAD! VDD_PAD! dn PJ=0.00041 m=1 $X=14104760 $Y=80300 $D=9
D2235 VDD_PAD! vdd! dn PJ=0.00041 m=1 $X=14107260 $Y=80300 $D=9
D2236 vdd! VDD_PAD! dn PJ=0.00041 m=1 $X=14109760 $Y=80300 $D=9
D2237 GND_PAD! VDD_PAD! dn PJ=0.00041 m=1 $X=14114760 $Y=80300 $D=9
D2238 VDD_PAD! vdd! dn PJ=0.00041 m=1 $X=14117260 $Y=80300 $D=9
D2239 vdd! VDD_PAD! dn PJ=0.00041 m=1 $X=14119760 $Y=80300 $D=9
D2240 GND_PAD! VDD_PAD! dn PJ=0.00041 m=1 $X=14124760 $Y=80300 $D=9
D2241 VDD_PAD! vdd! dn PJ=0.00041 m=1 $X=14127260 $Y=80300 $D=9
D2242 vdd! VDD_PAD! dn PJ=0.00041 m=1 $X=14129760 $Y=80300 $D=9
D2243 GND_PAD! VDD_PAD! dn PJ=0.00041 m=1 $X=14134760 $Y=80300 $D=9
D2244 VDD_PAD! vdd! dn PJ=0.00041 m=1 $X=14137260 $Y=80300 $D=9
D2245 vdd! VDD_PAD! dn PJ=0.00041 m=1 $X=14139760 $Y=80300 $D=9
D2246 GND_PAD! VDD_PAD! dn PJ=0.00041 m=1 $X=14144760 $Y=80300 $D=9
D2247 VDD_PAD! vdd! dn PJ=0.00041 m=1 $X=14147260 $Y=80300 $D=9
X2248 vdd! 534 534 pmos_a_CDNS_5887047866540 $T=12500 13207680 1 180 $X=11060 $Y=13207680
X2249 vdd! 584 584 pmos_a_CDNS_5887047866540 $T=14079860 13207680 1 180 $X=14078420 $Y=13207680
X2252 gnd! vdd! VDD_PAD $T=50000 180000 1 180 $X=-55000 $Y=-55000
X2253 gnd! vdd! VDD_PAD $T=3350000 180000 1 180 $X=3245000 $Y=-55000
X2254 gnd! vdd! VDD_PAD $T=3550000 180000 0 0 $X=3545000 $Y=-55000
X2255 gnd! vdd! VDD_PAD $T=7850000 180000 1 180 $X=7745000 $Y=-55000
X2256 gnd! vdd! VDD_PAD $T=10550000 180000 1 180 $X=10445000 $Y=-55000
X2257 gnd! vdd! VDD_PAD $T=10850000 180000 1 180 $X=10745000 $Y=-55000
X2258 gnd! vdd! VDD_PAD $T=14150000 180000 1 180 $X=14045000 $Y=-55000
X2261 181 78 nWE gnd! vdd! NWR 107 PADIN_WE $T=8920000 13542800 0 180 $X=8815000 $Y=13179780
X2262 191 154 193 gnd! vdd! BIT32 Bit_32 PADIN_WE $T=13860000 13542800 0 180 $X=13755000 $Y=13179780
X2263 194 154 196 gnd! vdd! BIT16 Bit_16 PADIN_WE $T=14120000 13542800 0 180 $X=14015000 $Y=13179780
X2264 gnd! vdd! gnd! vdd! PAD_Fill_160 $T=80000 13642800 1 0 $X=80000 $Y=13198800
X2265 gnd! vdd! gnd! vdd! PAD_Fill_160 $T=340000 13642800 1 0 $X=340000 $Y=13198800
X2266 gnd! vdd! gnd! vdd! PAD_Fill_160 $T=600000 13642800 1 0 $X=600000 $Y=13198800
X2267 gnd! vdd! gnd! vdd! PAD_Fill_160 $T=860000 13642800 1 0 $X=860000 $Y=13198800
X2268 gnd! vdd! gnd! vdd! PAD_Fill_160 $T=1380000 13642800 1 0 $X=1380000 $Y=13198800
X2269 gnd! vdd! gnd! vdd! PAD_Fill_160 $T=1640000 13642800 1 0 $X=1640000 $Y=13198800
X2270 gnd! vdd! gnd! vdd! PAD_Fill_160 $T=1900000 13642800 1 0 $X=1900000 $Y=13198800
X2271 gnd! vdd! gnd! vdd! PAD_Fill_160 $T=2160000 13642800 1 0 $X=2160000 $Y=13198800
X2272 gnd! vdd! gnd! vdd! PAD_Fill_160 $T=2420000 13642800 1 0 $X=2420000 $Y=13198800
X2273 gnd! vdd! gnd! vdd! PAD_Fill_160 $T=2680000 13642800 1 0 $X=2680000 $Y=13198800
X2274 gnd! vdd! gnd! vdd! PAD_Fill_160 $T=2940000 13642800 1 0 $X=2940000 $Y=13198800
X2275 gnd! vdd! gnd! vdd! PAD_Fill_160 $T=3200000 13642800 1 0 $X=3200000 $Y=13198800
X2276 gnd! vdd! gnd! vdd! PAD_Fill_160 $T=3460000 13642800 1 0 $X=3460000 $Y=13198800
X2277 gnd! vdd! gnd! vdd! PAD_Fill_160 $T=3720000 13642800 1 0 $X=3720000 $Y=13198800
X2278 gnd! vdd! gnd! vdd! PAD_Fill_160 $T=3980000 13642800 1 0 $X=3980000 $Y=13198800
X2279 gnd! vdd! gnd! vdd! PAD_Fill_160 $T=4240000 13642800 1 0 $X=4240000 $Y=13198800
X2280 gnd! vdd! gnd! vdd! PAD_Fill_160 $T=4500000 13642800 1 0 $X=4500000 $Y=13198800
X2281 gnd! vdd! gnd! vdd! PAD_Fill_160 $T=4760000 13642800 1 0 $X=4760000 $Y=13198800
X2282 gnd! vdd! gnd! vdd! PAD_Fill_160 $T=5280000 13642800 1 0 $X=5280000 $Y=13198800
X2283 gnd! vdd! gnd! vdd! PAD_Fill_160 $T=5540000 13642800 1 0 $X=5540000 $Y=13198800
X2284 gnd! vdd! gnd! vdd! PAD_Fill_160 $T=5800000 13642800 1 0 $X=5800000 $Y=13198800
X2285 gnd! vdd! gnd! vdd! PAD_Fill_160 $T=6060000 13642800 1 0 $X=6060000 $Y=13198800
X2286 gnd! vdd! gnd! vdd! PAD_Fill_160 $T=6320000 13642800 1 0 $X=6320000 $Y=13198800
X2287 gnd! vdd! gnd! vdd! PAD_Fill_160 $T=7780000 13642800 0 180 $X=7620000 $Y=13198800
X2288 gnd! vdd! gnd! vdd! PAD_Fill_160 $T=8040000 13642800 0 180 $X=7880000 $Y=13198800
X2289 gnd! vdd! gnd! vdd! PAD_Fill_160 $T=8300000 13642800 0 180 $X=8140000 $Y=13198800
X2290 gnd! vdd! gnd! vdd! PAD_Fill_160 $T=8560000 13642800 0 180 $X=8400000 $Y=13198800
X2291 gnd! vdd! gnd! vdd! PAD_Fill_160 $T=8820000 13642800 0 180 $X=8660000 $Y=13198800
X2292 gnd! vdd! gnd! vdd! PAD_Fill_160 $T=9080000 13642800 0 180 $X=8920000 $Y=13198800
X2293 gnd! vdd! gnd! vdd! PAD_Fill_160 $T=9340000 13642800 0 180 $X=9180000 $Y=13198800
X2294 gnd! vdd! gnd! vdd! PAD_Fill_160 $T=9860000 13642800 0 180 $X=9700000 $Y=13198800
X2295 gnd! vdd! gnd! vdd! PAD_Fill_160 $T=10120000 13642800 0 180 $X=9960000 $Y=13198800
X2296 gnd! vdd! gnd! vdd! PAD_Fill_160 $T=10380000 13642800 0 180 $X=10220000 $Y=13198800
X2297 gnd! vdd! gnd! vdd! PAD_Fill_160 $T=10640000 13642800 0 180 $X=10480000 $Y=13198800
X2298 gnd! vdd! gnd! vdd! PAD_Fill_160 $T=10900000 13642800 0 180 $X=10740000 $Y=13198800
X2299 gnd! vdd! gnd! vdd! PAD_Fill_160 $T=11160000 13642800 0 180 $X=11000000 $Y=13198800
X2300 gnd! vdd! gnd! vdd! PAD_Fill_160 $T=11420000 13642800 0 180 $X=11260000 $Y=13198800
X2301 gnd! vdd! gnd! vdd! PAD_Fill_160 $T=11680000 13642800 0 180 $X=11520000 $Y=13198800
X2302 gnd! vdd! gnd! vdd! PAD_Fill_160 $T=11940000 13642800 0 180 $X=11780000 $Y=13198800
X2303 gnd! vdd! gnd! vdd! PAD_Fill_160 $T=12200000 13642800 0 180 $X=12040000 $Y=13198800
X2304 gnd! vdd! gnd! vdd! PAD_Fill_160 $T=12460000 13642800 0 180 $X=12300000 $Y=13198800
X2305 gnd! vdd! gnd! vdd! PAD_Fill_160 $T=12720000 13642800 0 180 $X=12560000 $Y=13198800
X2306 gnd! vdd! gnd! vdd! PAD_Fill_160 $T=12980000 13642800 0 180 $X=12820000 $Y=13198800
X2307 gnd! vdd! gnd! vdd! PAD_Fill_160 $T=13500000 13642800 0 180 $X=13340000 $Y=13198800
X2308 gnd! vdd! gnd! vdd! PAD_Fill_160 $T=13760000 13642800 0 180 $X=13600000 $Y=13198800
X2309 gnd! vdd! gnd! vdd! PAD_Fill_160 $T=14020000 13642800 0 180 $X=13860000 $Y=13198800
X2310 GND_PAD! VDD_PAD! gnd! vdd! PAD_Fill_200 $T=2650000 80000 1 180 $X=2450000 $Y=-56000
X2311 GND_PAD! VDD_PAD! gnd! vdd! PAD_Fill_200 $T=2950000 80000 1 180 $X=2750000 $Y=-56000
X2312 GND_PAD! VDD_PAD! gnd! vdd! PAD_Fill_200 $T=3250000 80000 1 180 $X=3050000 $Y=-56000
X2313 GND_PAD! VDD_PAD! gnd! vdd! PAD_Fill_200 $T=3550000 80000 1 180 $X=3350000 $Y=-56000
X2314 GND_PAD! VDD_PAD! gnd! vdd! PAD_Fill_200 $T=6250000 80000 1 180 $X=6050000 $Y=-56000
X2315 GND_PAD! VDD_PAD! gnd! vdd! PAD_Fill_200 $T=6550000 80000 1 180 $X=6350000 $Y=-56000
X2316 GND_PAD! VDD_PAD! gnd! vdd! PAD_Fill_200 $T=6850000 80000 1 180 $X=6650000 $Y=-56000
X2317 GND_PAD! VDD_PAD! gnd! vdd! PAD_Fill_200 $T=7150000 80000 1 180 $X=6950000 $Y=-56000
X2318 GND_PAD! VDD_PAD! gnd! vdd! PAD_Fill_200 $T=7450000 80000 1 180 $X=7250000 $Y=-56000
X2319 GND_PAD! VDD_PAD! gnd! vdd! PAD_Fill_200 $T=7750000 80000 1 180 $X=7550000 $Y=-56000
X2320 GND_PAD! VDD_PAD! gnd! vdd! PAD_Fill_200 $T=10450000 80000 1 180 $X=10250000 $Y=-56000
X2321 GND_PAD! VDD_PAD! gnd! vdd! PAD_Fill_200 $T=10750000 80000 1 180 $X=10550000 $Y=-56000
X2322 GND_PAD! VDD_PAD! gnd! vdd! PAD_Fill_200 $T=11050000 80000 1 180 $X=10850000 $Y=-56000
X2323 GND_PAD! VDD_PAD! gnd! vdd! PAD_Fill_200 $T=11350000 80000 1 180 $X=11150000 $Y=-56000
X2324 GND_PAD! VDD_PAD! gnd! vdd! PAD_Fill_200 $T=14050000 80000 1 180 $X=13850000 $Y=-56000
X2325 Bit_32 gnd! 75 656 vdd! nOE_32 $T=3936560 518480 0 0 $X=3935740 $Y=511880
X2326 Bit_32 gnd! 75 655 vdd! nOE_32 $T=4236560 518480 0 0 $X=4235740 $Y=511880
X2327 Bit_32 gnd! 75 658 vdd! nOE_32 $T=4536560 518480 0 0 $X=4535740 $Y=511880
X2328 Bit_32 gnd! 75 657 vdd! nOE_32 $T=4836560 518480 0 0 $X=4835740 $Y=511880
X2329 Bit_32 gnd! 75 649 vdd! nOE_32 $T=5136560 518480 0 0 $X=5135740 $Y=511880
X2330 Bit_32 gnd! 75 660 vdd! nOE_32 $T=5436560 518480 0 0 $X=5435740 $Y=511880
X2331 Bit_32 gnd! 75 659 vdd! nOE_32 $T=5736560 518480 0 0 $X=5735740 $Y=511880
X2332 Bit_32 gnd! 75 652 vdd! nOE_32 $T=6036560 518480 0 0 $X=6035740 $Y=511880
X2333 Bit_32 gnd! 75 668 vdd! nOE_32 $T=11736560 518480 0 0 $X=11735740 $Y=511880
X2334 Bit_32 gnd! 75 667 vdd! nOE_32 $T=12036560 518480 0 0 $X=12035740 $Y=511880
X2335 Bit_32 gnd! 75 670 vdd! nOE_32 $T=12336560 518480 0 0 $X=12335740 $Y=511880
X2336 Bit_32 gnd! 75 669 vdd! nOE_32 $T=12636560 518480 0 0 $X=12635740 $Y=511880
X2337 Bit_32 gnd! 75 651 vdd! nOE_32 $T=12936560 518480 0 0 $X=12935740 $Y=511880
X2338 Bit_32 gnd! 75 672 vdd! nOE_32 $T=13236560 518480 0 0 $X=13235740 $Y=511880
X2339 Bit_32 gnd! 75 671 vdd! nOE_32 $T=13536560 518480 0 0 $X=13535740 $Y=511880
X2340 Bit_32 gnd! 75 654 vdd! nOE_32 $T=13836560 518480 0 0 $X=13835740 $Y=511880
X2341 Bit_16 Bit_32 280 87 317 318 DI_Bank<1> 319 DO_Bank<1> 4 vdd! gnd! 498 499 318 318 318 499 498 585 Select_Bit $T=290880 512020 0 0 $X=281500 $Y=500000
X2342 Bit_16 Bit_32 280 87 320 321 DI_Bank<2> 322 DO_Bank<2> 7 vdd! gnd! 500 501 321 321 321 501 500 586 Select_Bit $T=590880 512020 0 0 $X=581500 $Y=500000
X2343 Bit_16 Bit_32 280 87 323 324 DI_Bank<3> 325 DO_Bank<3> 9 vdd! gnd! 502 503 324 324 324 503 502 587 Select_Bit $T=890880 512020 0 0 $X=881500 $Y=500000
X2344 Bit_16 Bit_32 280 87 326 327 DI_Bank<4> 328 DO_Bank<4> 12 vdd! gnd! 504 505 327 327 327 505 504 588 Select_Bit $T=1190880 512020 0 0 $X=1181500 $Y=500000
X2345 Bit_16 Bit_32 280 87 329 330 DI_Bank<5> 331 DO_Bank<5> 15 vdd! gnd! 506 507 330 330 330 507 506 589 Select_Bit $T=1490880 512020 0 0 $X=1481500 $Y=500000
X2346 Bit_16 Bit_32 280 87 332 333 DI_Bank<6> 334 DO_Bank<6> 16 vdd! gnd! 508 509 333 333 333 509 508 590 Select_Bit $T=1790880 512020 0 0 $X=1781500 $Y=500000
X2347 Bit_16 Bit_32 280 87 335 336 DI_Bank<7> 337 DO_Bank<7> 22 vdd! gnd! 510 511 336 336 336 511 510 591 Select_Bit $T=2090880 512020 0 0 $X=2081500 $Y=500000
X2348 Bit_16 Bit_32 280 87 338 339 DI_Bank<8> 340 DO_Bank<8> 28 vdd! gnd! 512 513 339 339 339 513 512 592 Select_Bit $T=2390880 512020 0 0 $X=2381500 $Y=500000
X2349 Bit_16 Bit_32 280 87 341 DI_Bank<1> DI_Bank<17> 4 DO_Bank<17> 40 vdd! gnd! 87 514 593 550 550 514 594 550 Select_Bit $T=3890880 512020 0 0 $X=3881500 $Y=500000
X2350 Bit_16 Bit_32 280 87 342 DI_Bank<2> DI_Bank<18> 7 DO_Bank<18> 45 vdd! gnd! 87 515 595 551 551 515 596 551 Select_Bit $T=4190880 512020 0 0 $X=4181500 $Y=500000
X2351 Bit_16 Bit_32 280 87 343 DI_Bank<3> DI_Bank<19> 9 DO_Bank<19> 47 vdd! gnd! 87 516 597 552 552 516 598 552 Select_Bit $T=4490880 512020 0 0 $X=4481500 $Y=500000
X2352 Bit_16 Bit_32 280 87 344 DI_Bank<4> DI_Bank<20> 12 DO_Bank<20> 50 vdd! gnd! 87 517 599 553 553 517 600 553 Select_Bit $T=4790880 512020 0 0 $X=4781500 $Y=500000
X2353 Bit_16 Bit_32 280 87 345 DI_Bank<5> DI_Bank<21> 15 DO_Bank<21> 53 vdd! gnd! 87 518 601 554 554 518 602 554 Select_Bit $T=5090880 512020 0 0 $X=5081500 $Y=500000
X2354 Bit_16 Bit_32 280 87 346 DI_Bank<6> DI_Bank<22> 16 DO_Bank<22> 54 vdd! gnd! 87 519 603 555 555 519 604 555 Select_Bit $T=5390880 512020 0 0 $X=5381500 $Y=500000
X2355 Bit_16 Bit_32 280 87 347 DI_Bank<7> DI_Bank<23> 22 DO_Bank<23> 60 vdd! gnd! 87 520 605 556 556 520 606 556 Select_Bit $T=5690880 512020 0 0 $X=5681500 $Y=500000
X2356 Bit_16 Bit_32 280 87 348 DI_Bank<8> DI_Bank<24> 28 DO_Bank<24> 66 vdd! gnd! 87 521 607 557 557 521 608 557 Select_Bit $T=5990880 512020 0 0 $X=5981500 $Y=500000
X2357 Bit_16 Bit_32 280 87 349 DI_Bank<17> DI_Bank<9> 40 DO_Bank<9> 101 vdd! gnd! 522 280 609 609 564 610 522 564 Select_Bit $T=8090880 512020 0 0 $X=8081500 $Y=500000
X2358 Bit_16 Bit_32 280 87 350 DI_Bank<18> DI_Bank<10> 45 DO_Bank<10> 106 vdd! gnd! 523 280 611 611 565 612 523 565 Select_Bit $T=8390880 512020 0 0 $X=8381500 $Y=500000
X2359 Bit_16 Bit_32 280 87 351 DI_Bank<19> DI_Bank<11> 47 DO_Bank<11> 110 vdd! gnd! 524 280 613 613 566 614 524 566 Select_Bit $T=8690880 512020 0 0 $X=8681500 $Y=500000
X2360 Bit_16 Bit_32 280 87 352 DI_Bank<20> DI_Bank<12> 50 DO_Bank<12> 112 vdd! gnd! 525 280 615 615 567 616 525 567 Select_Bit $T=8990880 512020 0 0 $X=8981500 $Y=500000
X2361 Bit_16 Bit_32 280 87 353 DI_Bank<21> DI_Bank<13> 53 DO_Bank<13> 115 vdd! gnd! 526 280 617 617 568 618 526 568 Select_Bit $T=9290880 512020 0 0 $X=9281500 $Y=500000
X2362 Bit_16 Bit_32 280 87 354 DI_Bank<22> DI_Bank<14> 54 DO_Bank<14> 118 vdd! gnd! 527 280 619 619 569 620 527 569 Select_Bit $T=9590880 512020 0 0 $X=9581500 $Y=500000
X2363 Bit_16 Bit_32 280 87 355 DI_Bank<23> DI_Bank<15> 60 DO_Bank<15> 120 vdd! gnd! 528 280 621 621 570 622 528 570 Select_Bit $T=9890880 512020 0 0 $X=9881500 $Y=500000
X2364 Bit_16 Bit_32 280 87 356 DI_Bank<24> DI_Bank<16> 66 DO_Bank<16> 128 vdd! gnd! 529 280 623 623 571 624 529 571 Select_Bit $T=10190880 512020 0 0 $X=10181500 $Y=500000
X2365 Bit_16 Bit_32 280 87 357 DI_Bank<9> DI_Bank<25> 101 DO_Bank<25> gnd! vdd! gnd! 87 280 625 572 572 626 627 572 Select_Bit $T=11690880 512020 0 0 $X=11681500 $Y=500000
X2366 Bit_16 Bit_32 280 87 358 DI_Bank<10> DI_Bank<26> 106 DO_Bank<26> gnd! vdd! gnd! 87 280 628 573 573 629 630 573 Select_Bit $T=11990880 512020 0 0 $X=11981500 $Y=500000
X2367 Bit_16 Bit_32 280 87 359 DI_Bank<11> DI_Bank<27> 110 DO_Bank<27> gnd! vdd! gnd! 87 280 631 574 574 632 633 574 Select_Bit $T=12290880 512020 0 0 $X=12281500 $Y=500000
X2368 Bit_16 Bit_32 280 87 360 DI_Bank<12> DI_Bank<28> 112 DO_Bank<28> gnd! vdd! gnd! 87 280 634 575 575 635 636 575 Select_Bit $T=12590880 512020 0 0 $X=12581500 $Y=500000
X2369 Bit_16 Bit_32 280 87 361 DI_Bank<13> DI_Bank<29> 115 DO_Bank<29> gnd! vdd! gnd! 87 280 637 576 576 638 639 576 Select_Bit $T=12890880 512020 0 0 $X=12881500 $Y=500000
X2370 Bit_16 Bit_32 280 87 362 DI_Bank<14> DI_Bank<30> 118 DO_Bank<30> gnd! vdd! gnd! 87 280 640 577 577 641 642 577 Select_Bit $T=13190880 512020 0 0 $X=13181500 $Y=500000
X2371 Bit_16 Bit_32 280 87 363 DI_Bank<15> DI_Bank<31> 120 DO_Bank<31> gnd! vdd! gnd! 87 280 643 578 578 644 645 578 Select_Bit $T=13490880 512020 0 0 $X=13481500 $Y=500000
X2372 Bit_16 Bit_32 280 87 364 DI_Bank<16> DI_Bank<32> 128 DO_Bank<32> gnd! vdd! gnd! 87 280 646 579 579 647 648 579 Select_Bit $T=13790880 512020 0 0 $X=13781500 $Y=500000
X2373 gnd! vdd! Fill_Block_8Kx8 $T=3882880 524000 1 180 $X=3442680 $Y=523680
X2374 gnd! vdd! Fill_Block_8Kx8 $T=6966240 524000 1 180 $X=6526040 $Y=523680
X2375 gnd! vdd! Fill_Block_8Kx8 $T=8895680 524000 0 0 $X=8895320 $Y=523680
X2376 gnd! vdd! Fill_Block_8Kx8 $T=13740960 524000 0 0 $X=13740600 $Y=523680
X2377 80 GND_PAD! VDD_PAD! gnd! vdd! DIO5 329 331 75 PADIO $T=1450000 180000 0 0 $X=1445000 $Y=-55000
X2378 80 GND_PAD! VDD_PAD! gnd! vdd! DIO21 345 15 649 PADIO $T=5050000 180000 0 0 $X=5045000 $Y=-55000
X2379 80 GND_PAD! VDD_PAD! gnd! vdd! DIO13 353 53 650 PADIO $T=9250000 180000 0 0 $X=9245000 $Y=-55000
X2380 80 GND_PAD! VDD_PAD! gnd! vdd! DIO29 361 115 651 PADIO $T=12850000 180000 0 0 $X=12845000 $Y=-55000
X2381 GND_PAD! VDD_PAD! gnd! vdd! 80 DIO8 338 340 75 ICV_30 $T=2350000 80000 1 180 $X=2150000 $Y=-56000
X2382 GND_PAD! VDD_PAD! gnd! vdd! 80 DIO24 348 28 652 ICV_30 $T=5950000 80000 1 180 $X=5750000 $Y=-56000
X2383 GND_PAD! VDD_PAD! gnd! vdd! 80 DIO16 356 66 653 ICV_30 $T=10150000 80000 1 180 $X=9950000 $Y=-56000
X2384 GND_PAD! VDD_PAD! gnd! vdd! 80 DIO32 364 128 654 ICV_30 $T=13750000 80000 1 180 $X=13550000 $Y=-56000
X2385 gnd! vdd! GND_Core $T=600000 13542800 0 180 $X=495000 $Y=13198800
X2386 gnd! vdd! GND_Core $T=860000 13542800 0 180 $X=755000 $Y=13198800
X2387 gnd! vdd! GND_Core $T=2940000 13542800 0 180 $X=2835000 $Y=13198800
X2388 gnd! vdd! GND_Core $T=4500000 13542800 0 180 $X=4395000 $Y=13198800
X2389 gnd! vdd! GND_Core $T=4760000 13542800 0 180 $X=4655000 $Y=13198800
X2390 gnd! vdd! GND_Core $T=9700000 13542800 0 180 $X=9595000 $Y=13198800
X2391 gnd! vdd! GND_Core $T=9960000 13542800 0 180 $X=9855000 $Y=13198800
X2392 gnd! vdd! GND_Core $T=11520000 13542800 0 180 $X=11415000 $Y=13198800
X2393 gnd! vdd! GND_Core $T=13340000 13542800 0 180 $X=13235000 $Y=13198800
X2394 gnd! vdd! GND_Core $T=13600000 13542800 0 180 $X=13495000 $Y=13198800
X2395 gnd! vdd! PAD_Clamp_160 $T=1120000 13642800 1 0 $X=1120000 $Y=13198800
X2396 gnd! vdd! PAD_Clamp_160 $T=5020000 13642800 1 0 $X=5020000 $Y=13198800
X2397 gnd! vdd! PAD_Clamp_160 $T=9440000 13642800 1 0 $X=9440000 $Y=13198800
X2398 gnd! vdd! PAD_Clamp_160 $T=13080000 13642800 1 0 $X=13080000 $Y=13198800
X2399 vdd! gnd! VDD_Core $T=1380000 13542800 0 180 $X=1275000 $Y=13198800
X2400 vdd! gnd! VDD_Core $T=1640000 13542800 0 180 $X=1535000 $Y=13198800
X2401 vdd! gnd! VDD_Core $T=3200000 13542800 0 180 $X=3095000 $Y=13198800
X2402 vdd! gnd! VDD_Core $T=5020000 13542800 0 180 $X=4915000 $Y=13198800
X2403 vdd! gnd! VDD_Core $T=5280000 13542800 0 180 $X=5175000 $Y=13198800
X2404 vdd! gnd! VDD_Core $T=9180000 13542800 0 180 $X=9075000 $Y=13198800
X2405 vdd! gnd! VDD_Core $T=9440000 13542800 0 180 $X=9335000 $Y=13198800
X2406 vdd! gnd! VDD_Core $T=11260000 13542800 0 180 $X=11155000 $Y=13198800
X2407 vdd! gnd! VDD_Core $T=12820000 13542800 0 180 $X=12715000 $Y=13198800
X2408 vdd! gnd! VDD_Core $T=13080000 13542800 0 180 $X=12975000 $Y=13198800
X2409 GND_PAD! VDD_PAD! gnd! vdd! DIO2 80 DIO1 322 320 319 317 75 75 ICV_38 $T=250000 80000 1 180 $X=50000 $Y=-56000
X2410 GND_PAD! VDD_PAD! gnd! vdd! DIO4 80 DIO3 328 326 325 323 75 75 ICV_38 $T=850000 80000 1 180 $X=650000 $Y=-56000
X2411 GND_PAD! VDD_PAD! gnd! vdd! DIO7 80 DIO6 337 335 334 332 75 75 ICV_38 $T=1750000 80000 1 180 $X=1550000 $Y=-56000
X2412 GND_PAD! VDD_PAD! gnd! vdd! DIO18 80 DIO17 7 342 4 341 655 656 ICV_38 $T=3850000 80000 1 180 $X=3650000 $Y=-56000
X2413 GND_PAD! VDD_PAD! gnd! vdd! DIO20 80 DIO19 12 344 9 343 657 658 ICV_38 $T=4450000 80000 1 180 $X=4250000 $Y=-56000
X2414 GND_PAD! VDD_PAD! gnd! vdd! DIO23 80 DIO22 22 347 16 346 659 660 ICV_38 $T=5350000 80000 1 180 $X=5150000 $Y=-56000
X2415 GND_PAD! VDD_PAD! gnd! vdd! DIO10 80 DIO9 45 350 40 349 661 662 ICV_38 $T=8050000 80000 1 180 $X=7850000 $Y=-56000
X2416 GND_PAD! VDD_PAD! gnd! vdd! DIO12 80 DIO11 50 352 47 351 663 664 ICV_38 $T=8650000 80000 1 180 $X=8450000 $Y=-56000
X2417 GND_PAD! VDD_PAD! gnd! vdd! DIO15 80 DIO14 60 355 54 354 665 666 ICV_38 $T=9550000 80000 1 180 $X=9350000 $Y=-56000
X2418 GND_PAD! VDD_PAD! gnd! vdd! DIO26 80 DIO25 106 358 101 357 667 668 ICV_38 $T=11650000 80000 1 180 $X=11450000 $Y=-56000
X2419 GND_PAD! VDD_PAD! gnd! vdd! DIO28 80 DIO27 112 360 110 359 669 670 ICV_38 $T=12250000 80000 1 180 $X=12050000 $Y=-56000
X2420 GND_PAD! VDD_PAD! gnd! vdd! DIO31 80 DIO30 120 363 118 362 671 672 ICV_38 $T=13150000 80000 1 180 $X=12950000 $Y=-56000
X2421 gnd! vdd! ICV_39 $T=12860000 524000 0 0 $X=12859640 $Y=523680
X2422 VDD_PAD! vdd! gnd! GND_PAD! PAD_Clamp_200 $T=1450000 80000 1 180 $X=1250000 $Y=-56000
X2423 VDD_PAD! vdd! gnd! GND_PAD! PAD_Clamp_200 $T=5050000 80000 1 180 $X=4850000 $Y=-56000
X2424 VDD_PAD! vdd! gnd! GND_PAD! PAD_Clamp_200 $T=9250000 80000 1 180 $X=9050000 $Y=-56000
X2425 VDD_PAD! vdd! gnd! GND_PAD! PAD_Clamp_200 $T=12850000 80000 1 180 $X=12650000 $Y=-56000
X2426 78 gnd! vdd! A18 142 Bit_16 Bit_16 88 PADIN_Adress_Select $T=12200000 13542800 1 0 $X=12195000 $Y=13194180
X2427 78 gnd! vdd! A19 141 Bit_32 Bit_16 85 PADIN_Adress_Select $T=12460000 13542800 1 0 $X=12455000 $Y=13194180
X2428 gnd! vdd! ICV_83 $T=7133760 524000 0 0 $X=7133400 $Y=523680
X2429 gnd! vdd! ICV_83 $T=7133760 13198800 1 0 $X=7133400 $Y=13131600
X2430 gnd! vdd! ICV_83 $T=8895680 13198800 1 0 $X=8895320 $Y=13131600
X2431 gnd! vdd! ICV_83 $T=9336160 524000 0 0 $X=9335800 $Y=523680
X2432 gnd! vdd! ICV_83 $T=10657600 13198800 1 0 $X=10657240 $Y=13131600
X2433 gnd! vdd! ICV_83 $T=11098080 524000 0 0 $X=11097720 $Y=523680
X2434 gnd! vdd! ICV_83 $T=12419520 13198800 1 0 $X=12419160 $Y=13131600
X2435 23 18 25 365 679 680 gnd! vdd! RingPad_AND3 $T=2336160 13198800 0 0 $X=2335800 $Y=13198800
X2436 35 30 36 366 681 682 gnd! vdd! RingPad_AND3 $T=3636160 13198800 0 0 $X=3635800 $Y=13198800
X2437 56 57 61 367 683 684 gnd! vdd! RingPad_AND3 $T=5456160 13198800 0 0 $X=5455800 $Y=13198800
X2438 36 25 62 61 685 686 gnd! vdd! RingPad_AND3 $T=5717860 13198800 0 0 $X=5717500 $Y=13198800
X2439 93 94 104 368 687 688 gnd! vdd! RingPad_AND3 $T=7536160 13198800 0 0 $X=7535800 $Y=13198800
X2440 125 124 123 126 690 689 gnd! vdd! RingPad_AND3 $T=10202980 13198800 1 180 $X=10190660 $Y=13198800
X2441 312 127 124 312 691 692 gnd! vdd! RingPad_AND3 $T=10396160 13198800 0 0 $X=10395800 $Y=13198800
X2442 133 132 125 369 694 693 gnd! vdd! RingPad_AND3 $T=10723840 13198800 1 180 $X=10711520 $Y=13198800
X2443 142 141 126 370 696 695 gnd! vdd! RingPad_AND3 $T=12023840 13198800 1 180 $X=12011520 $Y=13198800
X2444 78 gnd! vdd! A0 18 Adr<0> PADIN_Adress $T=1900000 13542800 0 180 $X=1795000 $Y=13194180
X2445 78 gnd! vdd! A1 23 Adr<1> PADIN_Adress $T=2160000 13542800 0 180 $X=2055000 $Y=13194180
X2446 78 gnd! vdd! A2 365 Adr<2> PADIN_Adress $T=2320000 13542800 1 0 $X=2315000 $Y=13194180
X2447 78 gnd! vdd! A3 30 Adr<3> PADIN_Adress $T=2680000 13542800 0 180 $X=2575000 $Y=13194180
X2448 78 gnd! vdd! A4 35 Adr<4> PADIN_Adress $T=3460000 13542800 0 180 $X=3355000 $Y=13194180
X2449 78 gnd! vdd! A5 366 Adr<5> PADIN_Adress $T=3620000 13542800 1 0 $X=3615000 $Y=13194180
X2450 78 gnd! vdd! A6 57 Adr<6> PADIN_Adress $T=3980000 13542800 0 180 $X=3875000 $Y=13194180
X2451 78 gnd! vdd! A7 56 Adr<7> PADIN_Adress $T=4240000 13542800 0 180 $X=4135000 $Y=13194180
X2452 78 gnd! vdd! A8 367 Adr<8> PADIN_Adress $T=5440000 13542800 1 0 $X=5435000 $Y=13194180
X2453 78 gnd! vdd! A9 94 Adr<9> PADIN_Adress $T=5700000 13542800 1 0 $X=5695000 $Y=13194180
X2454 78 gnd! vdd! A10 93 Adr<10> PADIN_Adress $T=5960000 13542800 1 0 $X=5955000 $Y=13194180
X2455 78 gnd! vdd! A11 368 Adr<11> PADIN_Adress $T=7520000 13542800 1 0 $X=7515000 $Y=13194180
X2456 78 gnd! vdd! A12 127 83 PADIN_Adress $T=10220000 13542800 0 180 $X=10115000 $Y=13194180
X2457 78 gnd! vdd! A13 312 Adr<13> PADIN_Adress $T=10380000 13542800 1 0 $X=10375000 $Y=13194180
X2458 78 gnd! vdd! A14 369 Adr<14> PADIN_Adress $T=10740000 13542800 0 180 $X=10635000 $Y=13194180
X2459 78 gnd! vdd! A15 133 Adr<15> PADIN_Adress $T=10900000 13542800 1 0 $X=10895000 $Y=13194180
X2460 78 gnd! vdd! A16 132 Adr<16> PADIN_Adress $T=11680000 13542800 1 0 $X=11675000 $Y=13194180
X2461 78 gnd! vdd! A17 370 90 PADIN_Adress $T=12040000 13542800 0 180 $X=11935000 $Y=13194180
X2462 GND_PAD! VDD_PAD! gnd! vdd! GND_PAD $T=2750000 180000 1 180 $X=2645000 $Y=-55000
X2463 GND_PAD! VDD_PAD! gnd! vdd! GND_PAD $T=3050000 180000 1 180 $X=2945000 $Y=-55000
X2464 GND_PAD! VDD_PAD! gnd! vdd! GND_PAD $T=6350000 180000 1 180 $X=6245000 $Y=-55000
X2465 GND_PAD! VDD_PAD! gnd! vdd! GND_PAD $T=11150000 180000 1 180 $X=11045000 $Y=-55000
X2466 GND_PAD! VDD_PAD! gnd! vdd! GND_PAD $T=11450000 180000 1 180 $X=11345000 $Y=-55000
X2467 Bit_16 Bit_32 gnd! 75 662 vdd! nOE_16 $T=8136560 518480 0 0 $X=8135740 $Y=511840
X2468 Bit_16 Bit_32 gnd! 75 661 vdd! nOE_16 $T=8436560 518480 0 0 $X=8435740 $Y=511840
X2469 Bit_16 Bit_32 gnd! 75 664 vdd! nOE_16 $T=8736560 518480 0 0 $X=8735740 $Y=511840
X2470 Bit_16 Bit_32 gnd! 75 663 vdd! nOE_16 $T=9036560 518480 0 0 $X=9035740 $Y=511840
X2471 Bit_16 Bit_32 gnd! 75 650 vdd! nOE_16 $T=9336560 518480 0 0 $X=9335740 $Y=511840
X2472 Bit_16 Bit_32 gnd! 75 666 vdd! nOE_16 $T=9636560 518480 0 0 $X=9635740 $Y=511840
X2473 Bit_16 Bit_32 gnd! 75 665 vdd! nOE_16 $T=9936560 518480 0 0 $X=9935740 $Y=511840
X2474 Bit_16 Bit_32 gnd! 75 653 vdd! nOE_16 $T=10236560 518480 0 0 $X=10235740 $Y=511840
X2475 gnd! vdd! OEN 107 103 nOE_Core 76 PADIN_OE $T=8660000 13542800 0 180 $X=8555000 $Y=13177380
X2476 181 123 62 97 78 gnd! vdd! CEN 104 103 PADIN_CE $T=8400000 13542800 0 180 $X=8295000 $Y=13167780
X2477 gnd! vdd! Test 1 92 PADIN_CS $T=80000 13542800 0 180 $X=-25000 $Y=13177380
X2478 gnd! vdd! 252 1 371 PADIN_CS $T=340000 13542800 0 180 $X=235000 $Y=13177380
X2479 gnd! vdd! MODE 1 68 PADIN_CS $T=1020000 13542800 1 0 $X=1015000 $Y=13177380
X2480 gnd! vdd! A20 68 70 PADIN_CS $T=6320000 13542800 0 180 $X=6215000 $Y=13177380
X2481 gnd! vdd! CS1 68 306 PADIN_CS $T=6480000 13542800 1 0 $X=6475000 $Y=13177380
X2482 gnd! vdd! CS2 68 311 PADIN_CS $T=7880000 13542800 0 180 $X=7775000 $Y=13177380
X2483 gnd! vdd! A21 68 99 PADIN_CS $T=8140000 13542800 0 180 $X=8035000 $Y=13177380
X2486 306 70 98 gnd! vdd! 697 RingPad_EOR $T=6550220 13211280 1 0 $X=6545420 $Y=13198800
X2487 311 99 563 gnd! vdd! 698 RingPad_EOR $T=7809780 13211280 0 180 $X=7800660 $Y=13198800
X2488 vdd! gnd! VDD_Core_PAD $T=7250000 180000 1 180 $X=7145000 $Y=-55000
X2489 vdd! gnd! VDD_Core_PAD $T=7450000 180000 0 0 $X=7445000 $Y=-55000
X2490 76 75 vdd! gnd! RingPad_Buffer $T=7044660 555340 0 180 $X=7014300 $Y=551380
X2491 78 nCE vdd! gnd! RingPad_Buffer $T=7057060 13167460 1 180 $X=7026700 $Y=13166940
X2492 83 Adr<12> vdd! gnd! RingPad_Buffer $T=7087820 13167460 1 180 $X=7057460 $Y=13166940
X2493 Adr<19> 280 vdd! gnd! RingPad_Buffer $T=7095320 574560 0 180 $X=7064960 $Y=570600
X2494 85 Adr<19> vdd! gnd! RingPad_Buffer $T=7095340 13148240 1 180 $X=7064980 $Y=13147720
X2495 nWE 80 vdd! gnd! RingPad_Buffer $T=7072260 555340 1 0 $X=7072260 $Y=551380
X2496 88 Adr<18> vdd! gnd! RingPad_Buffer $T=7088220 13167460 0 0 $X=7088220 $Y=13166940
X2497 90 Adr<17> vdd! gnd! RingPad_Buffer $T=7095740 13148240 0 0 $X=7095740 $Y=13147720
X2498 Adr<18> 87 vdd! gnd! RingPad_Buffer $T=7095840 574560 1 0 $X=7095840 $Y=570600
X2499 vdd! gnd! Fill_Dec_X512 $T=7050040 589960 0 180 $X=6966240 $Y=523680
X2500 vdd! gnd! Fill_Dec_X512 $T=7050040 13132840 1 180 $X=6966240 $Y=13133240
X2501 vdd! gnd! Fill_Dec_X512 $T=7049960 589960 1 0 $X=7050000 $Y=523680
X2502 vdd! gnd! Fill_Dec_X512 $T=7049960 13132840 0 0 $X=7050000 $Y=13133240
X2503 gnd! GND_PAD! vdd! GND_Core_PAD $T=6650000 180000 1 180 $X=6545000 $Y=-55000
X2504 gnd! GND_PAD! vdd! GND_Core_PAD $T=6950000 180000 1 180 $X=6845000 $Y=-55000
X2505 gnd! vdd! 92 Usub Usub_7V $T=6505000 13492800 0 180 $X=6580000 $Y=13172580
X2506 gnd! vdd! ICV_166 $T=6085280 524000 1 180 $X=5645080 $Y=523680
X2507 gnd! vdd! ICV_167 $T=359040 524000 1 180 $X=-81160 $Y=523680
X2508 gnd! vdd! ICV_167 $T=359040 13198800 0 180 $X=-81160 $Y=13131600
X2509 gnd! vdd! ICV_167 $T=2120960 524000 1 180 $X=1680760 $Y=523680
X2510 gnd! vdd! ICV_167 $T=2120960 13198800 0 180 $X=1680760 $Y=13131600
X2511 gnd! vdd! ICV_167 $T=3882880 13198800 0 180 $X=3442680 $Y=13131600
X2512 gnd! vdd! ICV_167 $T=4323360 524000 1 180 $X=3883160 $Y=523680
X2513 gnd! vdd! ICV_167 $T=5644800 13198800 0 180 $X=5204600 $Y=13131600
.ENDS
***************************************
